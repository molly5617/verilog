//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

//added by CIC
`timescale 1ns/1ps
`celldefine
module ANTENNATH ( A );
    input A ;
endmodule
`endcelldefine

`timescale 1ns/1ps
`celldefine
module ACCSHCINX2TH ( CO0, CO1, A, B, CI0N, CI1N);
output CO0, CO1;
input A, B, CI0N, CI1N;
  not I0 (cin1, CI1N);
  not I1 (cin0, CI0N);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci0, A, cin0);
  and I4 (b_and_ci0, B, cin0);
  or  I5 (CO0, a_and_b, a_and_ci0, b_and_ci0);
  and I6 (a_and_ci1, A, cin1);
  and I7 (b_and_ci1, B, cin1);
  or  I8 (CO1, a_and_b, a_and_ci1, b_and_ci1);
  specify
    specparam

      tplh$A$CO0  = 1.0,
      tphl$A$CO0  = 1.0,
      tplh$A$CO1  = 1.0,
      tphl$A$CO1  = 1.0,
      tplh$B$CO0  = 1.0,
      tphl$B$CO0  = 1.0,
      tplh$B$CO1  = 1.0,
      tphl$B$CO1  = 1.0,
      tplh$CI0N$CO0  = 1.0,
      tphl$CI0N$CO0  = 1.0,
      tplh$CI0N$CO1  = 1.0,
      tphl$CI0N$CO1  = 1.0,
      tplh$CI1N$CO0  = 1.0,
      tphl$CI1N$CO0  = 1.0,
      tplh$CI1N$CO1  = 1.0,
      tphl$CI1N$CO1  = 1.0;


    if (A == 1'b1 && B == 1'b0 )
       (CI1N *> CO1) = (tplh$CI1N$CO1, tphl$CI1N$CO1); 
    if (A == 1'b0 && B == 1'b1 )
       (CI1N *> CO1) = (tplh$CI1N$CO1, tphl$CI1N$CO1); 
    if (A == 1'b1 && CI1N == 1'b1 )
       (B *> CO1) = (tplh$B$CO1, tphl$B$CO1); 
    if (A == 1'b0 && CI1N == 1'b0 )
       (B *> CO1) = (tplh$B$CO1, tphl$B$CO1); 
    if (B == 1'b1 && CI1N == 1'b1 )
       (A *> CO1) = (tplh$A$CO1, tphl$A$CO1); 
    if (B == 1'b0 && CI1N == 1'b0 )
       (A *> CO1) = (tplh$A$CO1, tphl$A$CO1); 
    if (A == 1'b1 && CI0N == 1'b1 )
       (B *> CO0) = (tplh$B$CO0, tphl$B$CO0); 
    if (A == 1'b0 && CI0N == 1'b0 )
       (B *> CO0) = (tplh$B$CO0, tphl$B$CO0); 
    if (B == 1'b1 && CI0N == 1'b1 )
       (A *> CO0) = (tplh$A$CO0, tphl$A$CO0); 
    if (B == 1'b0 && CI0N == 1'b0 )
       (A *> CO0) = (tplh$A$CO0, tphl$A$CO0); 
    if (A == 1'b1 && B == 1'b0 )
       (CI0N *> CO0) = (tplh$CI0N$CO0, tphl$CI0N$CO0); 
    if (A == 1'b0 && B == 1'b1 )
       (CI0N *> CO0) = (tplh$CI0N$CO0, tphl$CI0N$CO0);

  endspecify
endmodule // ACCSHCINX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ACCSHCINX4TH ( CO0, CO1, A, B, CI0N, CI1N);
output CO0, CO1;
input A, B, CI0N, CI1N;
  not I0 (cin1, CI1N);
  not I1 (cin0, CI0N);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci0, A, cin0);
  and I4 (b_and_ci0, B, cin0);
  or  I5 (CO0, a_and_b, a_and_ci0, b_and_ci0);
  and I6 (a_and_ci1, A, cin1);
  and I7 (b_and_ci1, B, cin1);
  or  I8 (CO1, a_and_b, a_and_ci1, b_and_ci1);
  specify
    specparam

      tplh$A$CO0  = 1.0,
      tphl$A$CO0  = 1.0,
      tplh$A$CO1  = 1.0,
      tphl$A$CO1  = 1.0,
      tplh$B$CO0  = 1.0,
      tphl$B$CO0  = 1.0,
      tplh$B$CO1  = 1.0,
      tphl$B$CO1  = 1.0,
      tplh$CI0N$CO0  = 1.0,
      tphl$CI0N$CO0  = 1.0,
      tplh$CI0N$CO1  = 1.0,
      tphl$CI0N$CO1  = 1.0,
      tplh$CI1N$CO0  = 1.0,
      tphl$CI1N$CO0  = 1.0,
      tplh$CI1N$CO1  = 1.0,
      tphl$CI1N$CO1  = 1.0;


    if (A == 1'b1 && B == 1'b0 )
       (CI1N *> CO1) = (tplh$CI1N$CO1, tphl$CI1N$CO1); 
    if (A == 1'b0 && B == 1'b1 )
       (CI1N *> CO1) = (tplh$CI1N$CO1, tphl$CI1N$CO1); 
    if (A == 1'b1 && CI1N == 1'b1 )
       (B *> CO1) = (tplh$B$CO1, tphl$B$CO1); 
    if (A == 1'b0 && CI1N == 1'b0 )
       (B *> CO1) = (tplh$B$CO1, tphl$B$CO1); 
    if (B == 1'b1 && CI1N == 1'b1 )
       (A *> CO1) = (tplh$A$CO1, tphl$A$CO1); 
    if (B == 1'b0 && CI1N == 1'b0 )
       (A *> CO1) = (tplh$A$CO1, tphl$A$CO1); 
    if (A == 1'b1 && CI0N == 1'b1 )
       (B *> CO0) = (tplh$B$CO0, tphl$B$CO0); 
    if (A == 1'b0 && CI0N == 1'b0 )
       (B *> CO0) = (tplh$B$CO0, tphl$B$CO0); 
    if (B == 1'b1 && CI0N == 1'b1 )
       (A *> CO0) = (tplh$A$CO0, tphl$A$CO0); 
    if (B == 1'b0 && CI0N == 1'b0 )
       (A *> CO0) = (tplh$A$CO0, tphl$A$CO0); 
    if (A == 1'b1 && B == 1'b0 )
       (CI0N *> CO0) = (tplh$CI0N$CO0, tphl$CI0N$CO0); 
    if (A == 1'b0 && B == 1'b1 )
       (CI0N *> CO0) = (tplh$CI0N$CO0, tphl$CI0N$CO0);

  endspecify
endmodule // ACCSHCINX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ACCSHCONX2TH ( CO0N, CO1N, A, B, CI0, CI1);
output CO0N, CO1N;
input A, B, CI0, CI1;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci0, A, CI0);
  and I2 (b_and_ci0, B, CI0);
  or  I3 (cout0, a_and_b, a_and_ci0, b_and_ci0);
  and I4 (a_and_ci1, A, CI1);
  and I5 (b_and_ci1, B, CI1);
  or  I6 (cout1, a_and_b, a_and_ci1, b_and_ci1);
  not I7 (CO1N, cout1);
  not I8 (CO0N, cout0);
  specify
    specparam

      tplh$A$CO0N  = 1.0,
      tphl$A$CO0N  = 1.0,
      tplh$A$CO1N  = 1.0,
      tphl$A$CO1N  = 1.0,
      tplh$B$CO0N  = 1.0,
      tphl$B$CO0N  = 1.0,
      tplh$B$CO1N  = 1.0,
      tphl$B$CO1N  = 1.0,
      tplh$CI0$CO0N  = 1.0,
      tphl$CI0$CO0N  = 1.0,
      tplh$CI0$CO1N  = 1.0,
      tphl$CI0$CO1N  = 1.0,
      tplh$CI1$CO0N  = 1.0,
      tphl$CI1$CO0N  = 1.0,
      tplh$CI1$CO1N  = 1.0,
      tphl$CI1$CO1N  = 1.0;


    if (B == 1'b1 && CI0 == 1'b0 )
       (A *> CO0N) = (tplh$A$CO0N, tphl$A$CO0N); 
    if (B == 1'b0 && CI0 == 1'b1 )
       (A *> CO0N) = (tplh$A$CO0N, tphl$A$CO0N); 
    if (A == 1'b1 && B == 1'b0 )
       (CI0 *> CO0N) = (tplh$CI0$CO0N, tphl$CI0$CO0N); 
    if (A == 1'b0 && B == 1'b1 )
       (CI0 *> CO0N) = (tplh$CI0$CO0N, tphl$CI0$CO0N); 
    if (A == 1'b1 && CI0 == 1'b0 )
       (B *> CO0N) = (tplh$B$CO0N, tphl$B$CO0N); 
    if (A == 1'b0 && CI0 == 1'b1 )
       (B *> CO0N) = (tplh$B$CO0N, tphl$B$CO0N); 
    if (B == 1'b1 && CI1 == 1'b0 )
       (A *> CO1N) = (tplh$A$CO1N, tphl$A$CO1N); 
    if (B == 1'b0 && CI1 == 1'b1 )
       (A *> CO1N) = (tplh$A$CO1N, tphl$A$CO1N); 
    if (A == 1'b1 && CI1 == 1'b0 )
       (B *> CO1N) = (tplh$B$CO1N, tphl$B$CO1N); 
    if (A == 1'b0 && CI1 == 1'b1 )
       (B *> CO1N) = (tplh$B$CO1N, tphl$B$CO1N); 
    if (A == 1'b1 && B == 1'b0 )
       (CI1 *> CO1N) = (tplh$CI1$CO1N, tphl$CI1$CO1N); 
    if (A == 1'b0 && B == 1'b1 )
       (CI1 *> CO1N) = (tplh$CI1$CO1N, tphl$CI1$CO1N);

  endspecify
endmodule // ACCSHCONX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ACCSHCONX4TH ( CO0N, CO1N, A, B, CI0, CI1);
output CO0N, CO1N;
input A, B, CI0, CI1;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci0, A, CI0);
  and I2 (b_and_ci0, B, CI0);
  or  I3 (cout0, a_and_b, a_and_ci0, b_and_ci0);
  and I4 (a_and_ci1, A, CI1);
  and I5 (b_and_ci1, B, CI1);
  or  I6 (cout1, a_and_b, a_and_ci1, b_and_ci1);
  not I7 (CO1N, cout1);
  not I8 (CO0N, cout0);
  specify
    specparam

      tplh$A$CO0N  = 1.0,
      tphl$A$CO0N  = 1.0,
      tplh$A$CO1N  = 1.0,
      tphl$A$CO1N  = 1.0,
      tplh$B$CO0N  = 1.0,
      tphl$B$CO0N  = 1.0,
      tplh$B$CO1N  = 1.0,
      tphl$B$CO1N  = 1.0,
      tplh$CI0$CO0N  = 1.0,
      tphl$CI0$CO0N  = 1.0,
      tplh$CI0$CO1N  = 1.0,
      tphl$CI0$CO1N  = 1.0,
      tplh$CI1$CO0N  = 1.0,
      tphl$CI1$CO0N  = 1.0,
      tplh$CI1$CO1N  = 1.0,
      tphl$CI1$CO1N  = 1.0;


    if (B == 1'b1 && CI0 == 1'b0 )
       (A *> CO0N) = (tplh$A$CO0N, tphl$A$CO0N); 
    if (B == 1'b0 && CI0 == 1'b1 )
       (A *> CO0N) = (tplh$A$CO0N, tphl$A$CO0N); 
    if (A == 1'b1 && B == 1'b0 )
       (CI0 *> CO0N) = (tplh$CI0$CO0N, tphl$CI0$CO0N); 
    if (A == 1'b0 && B == 1'b1 )
       (CI0 *> CO0N) = (tplh$CI0$CO0N, tphl$CI0$CO0N); 
    if (A == 1'b1 && CI0 == 1'b0 )
       (B *> CO0N) = (tplh$B$CO0N, tphl$B$CO0N); 
    if (A == 1'b0 && CI0 == 1'b1 )
       (B *> CO0N) = (tplh$B$CO0N, tphl$B$CO0N); 
    if (B == 1'b1 && CI1 == 1'b0 )
       (A *> CO1N) = (tplh$A$CO1N, tphl$A$CO1N); 
    if (B == 1'b0 && CI1 == 1'b1 )
       (A *> CO1N) = (tplh$A$CO1N, tphl$A$CO1N); 
    if (A == 1'b1 && CI1 == 1'b0 )
       (B *> CO1N) = (tplh$B$CO1N, tphl$B$CO1N); 
    if (A == 1'b0 && CI1 == 1'b1 )
       (B *> CO1N) = (tplh$B$CO1N, tphl$B$CO1N); 
    if (A == 1'b1 && B == 1'b0 )
       (CI1 *> CO1N) = (tplh$CI1$CO1N, tphl$CI1$CO1N); 
    if (A == 1'b0 && B == 1'b1 )
       (CI1 *> CO1N) = (tplh$CI1$CO1N, tphl$CI1$CO1N);

  endspecify
endmodule // ACCSHCONX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ACCSIHCONX2TH ( CO0N, CO1N, A, B);
output CO0N, CO1N;
input A, B;
  and I0 (CO0, A, B);
  or  I1 (CO1, A, B);
  not I2 (CO0N, CO0);
  not I3 (CO1N, CO1);
  specify
    specparam

      tplh$A$CO0N  = 1.0,
      tphl$A$CO0N  = 1.0,
      tplh$A$CO1N  = 1.0,
      tphl$A$CO1N  = 1.0,
      tplh$B$CO0N  = 1.0,
      tphl$B$CO0N  = 1.0,
      tplh$B$CO1N  = 1.0,
      tphl$B$CO1N  = 1.0;


	(A  *> CO0N)  = (tplh$A$CO0N,   tphl$A$CO0N);
	(B  *> CO0N)  = (tplh$B$CO0N,   tphl$B$CO0N);
	(A  *> CO1N)  = (tplh$A$CO1N,   tphl$A$CO1N);
	(B  *> CO1N)  = (tplh$B$CO1N,   tphl$B$CO1N);

  endspecify
endmodule // ACCSIHCONX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ACCSIHCONX4TH ( CO0N, CO1N, A, B);
output CO0N, CO1N;
input A, B;
  and I0 (CO0, A, B);
  or  I1 (CO1, A, B);
  not I2 (CO0N, CO0);
  not I3 (CO1N, CO1);
  specify
    specparam

      tplh$A$CO0N  = 1.0,
      tphl$A$CO0N  = 1.0,
      tplh$A$CO1N  = 1.0,
      tphl$A$CO1N  = 1.0,
      tplh$B$CO0N  = 1.0,
      tphl$B$CO0N  = 1.0,
      tplh$B$CO1N  = 1.0,
      tphl$B$CO1N  = 1.0;


	(A  *> CO0N)  = (tplh$A$CO0N,   tphl$A$CO0N);
	(B  *> CO0N)  = (tplh$B$CO0N,   tphl$B$CO0N);
	(A  *> CO1N)  = (tplh$A$CO1N,   tphl$A$CO1N);
	(B  *> CO1N)  = (tplh$B$CO1N,   tphl$B$CO1N);

  endspecify
endmodule // ACCSIHCONX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ACHCINX2TH ( CO, A, B, CIN);
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or  I4 (CO, a_and_b, a_and_ci, b_and_ci);   
  specify
    specparam

      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CIN$CO  = 1.0,
      tphl$CIN$CO  = 1.0;


    if (A == 1'b1 && B == 1'b0 )
       (CIN *> CO) = (tplh$CIN$CO, tphl$CIN$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CIN *> CO) = (tplh$CIN$CO, tphl$CIN$CO); 
    if (B == 1'b1 && CIN == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CIN == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CIN == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CIN == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO);

  endspecify
endmodule // ACHCINX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ACHCINX4TH ( CO, A, B, CIN);
output CO;
input A, B, CIN;
  and I0 (a_and_b, A, B);
  not I1 (ci, CIN);
  and I2 (a_and_ci, A, ci);
  and I3 (b_and_ci, B, ci);
  or  I4 (CO, a_and_b, a_and_ci, b_and_ci);   
  specify
    specparam

      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CIN$CO  = 1.0,
      tphl$CIN$CO  = 1.0;


    if (A == 1'b1 && B == 1'b0 )
       (CIN *> CO) = (tplh$CIN$CO, tphl$CIN$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CIN *> CO) = (tplh$CIN$CO, tphl$CIN$CO); 
    if (B == 1'b1 && CIN == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CIN == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CIN == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CIN == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO);

  endspecify
endmodule // ACHCINX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ACHCONX2TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or  I3 (cout, a_and_b, a_and_ci, b_and_ci);   
  not I4 (CON, cout);
  specify
    specparam

      tplh$A$CON  = 1.0,
      tphl$A$CON  = 1.0,
      tplh$B$CON  = 1.0,
      tphl$B$CON  = 1.0,
      tplh$CI$CON  = 1.0,
      tphl$CI$CON  = 1.0;


    if (B == 1'b1 && CI == 1'b0 )
       (A *> CON) = (tplh$A$CON, tphl$A$CON); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CON) = (tplh$A$CON, tphl$A$CON); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CON) = (tplh$B$CON, tphl$B$CON); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CON) = (tplh$B$CON, tphl$B$CON); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CON) = (tplh$CI$CON, tphl$CI$CON); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CON) = (tplh$CI$CON, tphl$CI$CON);

  endspecify
endmodule // ACHCONX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ACHCONX4TH ( CON, A, B, CI);
output CON;
input A, B, CI;
  and I0 (a_and_b, A, B);
  and I1 (a_and_ci, A, CI);
  and I2 (b_and_ci, B, CI);
  or  I3 (cout, a_and_b, a_and_ci, b_and_ci);   
  not I4 (CON, cout);
  specify
    specparam

      tplh$A$CON  = 1.0,
      tphl$A$CON  = 1.0,
      tplh$B$CON  = 1.0,
      tphl$B$CON  = 1.0,
      tplh$CI$CON  = 1.0,
      tphl$CI$CON  = 1.0;


    if (B == 1'b1 && CI == 1'b0 )
       (A *> CON) = (tplh$A$CON, tphl$A$CON); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CON) = (tplh$A$CON, tphl$A$CON); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CON) = (tplh$B$CON, tphl$B$CON); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CON) = (tplh$B$CON, tphl$B$CON); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CON) = (tplh$CI$CON, tphl$CI$CON); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CON) = (tplh$CI$CON, tphl$CI$CON);

  endspecify
endmodule // ACHCONX4TH
`endcelldefine
//$Id: cmpr.genpp,v 1.8 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CMPR42X1TH (S, CO, ICO, A, B, C, D, ICI);
output S, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or  I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor I7 (S, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or  I11 (CO, t5, t6, t7);
  specify
    // delay parameters
    specparam
      tplh$A$S = 1.0,
      tphl$A$S = 1.0,
      tplh$B$S = 1.0,
      tphl$B$S = 1.0,
      tplh$C$S = 1.0,
      tphl$C$S = 1.0,
      tplh$D$S = 1.0,
      tphl$D$S = 1.0,
      tplh$ICI$S = 1.0,
      tphl$ICI$S = 1.0,
      tplh$A$CO = 1.0,
      tphl$A$CO = 1.0,
      tplh$B$CO = 1.0,
      tphl$B$CO = 1.0,
      tplh$C$CO = 1.0,
      tphl$C$CO = 1.0,
      tplh$D$CO = 1.0,
      tphl$D$CO = 1.0,
      tplh$ICI$CO = 1.0,
      tphl$ICI$CO = 1.0,
      tplh$A$ICO = 1.0,
      tphl$A$ICO = 1.0,
      tplh$B$ICO = 1.0,
      tphl$B$ICO = 1.0,
      tplh$C$ICO = 1.0,
      tphl$C$ICO = 1.0,
      tplh$D$ICO = 1.0,
      tphl$D$ICO = 1.0,
      tplh$ICI$ICO = 1.0,
      tphl$ICI$ICO = 1.0;
    // path delays
     if (B == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) 
	(A *> S) = (tplh$A$S, tphl$A$S);
     if (!(B == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) )
	(A *> S) = (tplh$A$S, tphl$A$S);
     if (A == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) 
	(B *> S) = (tplh$B$S, tphl$B$S);
     if (!(A == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) )
	(B *> S) = (tplh$B$S, tphl$B$S);
     if (A == 1'b1 ^ B == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1)
	(C *> S) = (tplh$C$S, tphl$C$S);
     if (!(A == 1'b1 ^ B == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1))
	(C *> S) = (tplh$C$S, tphl$C$S);
     if (A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ ICI == 1'b1)
	(D *> S) = (tplh$D$S, tphl$D$S);
     if (!(A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ ICI == 1'b1))
	(D *> S) = (tplh$D$S, tphl$D$S);
     if (A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ D == 1'b1)
	(ICI *> S) = (tplh$ICI$S, tphl$ICI$S);
     if (!(A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ D == 1'b1))
	(ICI *> S) = (tplh$ICI$S, tphl$ICI$S);
    if (B == 1'b1 && C == 1'b0 )
       (A *> ICO) = (tplh$A$ICO, tphl$A$ICO); 
    if (B == 1'b0 && C == 1'b1 )
       (A *> ICO) = (tplh$A$ICO, tphl$A$ICO); 
    if (A == 1'b1 && C == 1'b0 )
       (B *> ICO) = (tplh$B$ICO, tphl$B$ICO); 
    if (A == 1'b0 && C == 1'b1 )
       (B *> ICO) = (tplh$B$ICO, tphl$B$ICO); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> ICO) = (tplh$C$ICO, tphl$C$ICO); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> ICO) = (tplh$C$ICO, tphl$C$ICO); 
    if (B == 1'b0 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b0 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && B == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO);
 
  endspecify

endmodule // CMPR42X1TH
`endcelldefine
//$Id: cmpr.genpp,v 1.8 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CMPR42X2TH (S, CO, ICO, A, B, C, D, ICI);
output S, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or  I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor I7 (S, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or  I11 (CO, t5, t6, t7);
  specify
    // delay parameters
    specparam
      tplh$A$S = 1.0,
      tphl$A$S = 1.0,
      tplh$B$S = 1.0,
      tphl$B$S = 1.0,
      tplh$C$S = 1.0,
      tphl$C$S = 1.0,
      tplh$D$S = 1.0,
      tphl$D$S = 1.0,
      tplh$ICI$S = 1.0,
      tphl$ICI$S = 1.0,
      tplh$A$CO = 1.0,
      tphl$A$CO = 1.0,
      tplh$B$CO = 1.0,
      tphl$B$CO = 1.0,
      tplh$C$CO = 1.0,
      tphl$C$CO = 1.0,
      tplh$D$CO = 1.0,
      tphl$D$CO = 1.0,
      tplh$ICI$CO = 1.0,
      tphl$ICI$CO = 1.0,
      tplh$A$ICO = 1.0,
      tphl$A$ICO = 1.0,
      tplh$B$ICO = 1.0,
      tphl$B$ICO = 1.0,
      tplh$C$ICO = 1.0,
      tphl$C$ICO = 1.0,
      tplh$D$ICO = 1.0,
      tphl$D$ICO = 1.0,
      tplh$ICI$ICO = 1.0,
      tphl$ICI$ICO = 1.0;
    // path delays
     if (B == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) 
	(A *> S) = (tplh$A$S, tphl$A$S);
     if (!(B == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) )
	(A *> S) = (tplh$A$S, tphl$A$S);
     if (A == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) 
	(B *> S) = (tplh$B$S, tphl$B$S);
     if (!(A == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) )
	(B *> S) = (tplh$B$S, tphl$B$S);
     if (A == 1'b1 ^ B == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1)
	(C *> S) = (tplh$C$S, tphl$C$S);
     if (!(A == 1'b1 ^ B == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1))
	(C *> S) = (tplh$C$S, tphl$C$S);
     if (A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ ICI == 1'b1)
	(D *> S) = (tplh$D$S, tphl$D$S);
     if (!(A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ ICI == 1'b1))
	(D *> S) = (tplh$D$S, tphl$D$S);
     if (A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ D == 1'b1)
	(ICI *> S) = (tplh$ICI$S, tphl$ICI$S);
     if (!(A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ D == 1'b1))
	(ICI *> S) = (tplh$ICI$S, tphl$ICI$S);
    if (B == 1'b1 && C == 1'b0 )
       (A *> ICO) = (tplh$A$ICO, tphl$A$ICO); 
    if (B == 1'b0 && C == 1'b1 )
       (A *> ICO) = (tplh$A$ICO, tphl$A$ICO); 
    if (A == 1'b1 && C == 1'b0 )
       (B *> ICO) = (tplh$B$ICO, tphl$B$ICO); 
    if (A == 1'b0 && C == 1'b1 )
       (B *> ICO) = (tplh$B$ICO, tphl$B$ICO); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> ICO) = (tplh$C$ICO, tphl$C$ICO); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> ICO) = (tplh$C$ICO, tphl$C$ICO); 
    if (B == 1'b0 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b0 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && B == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO);
 
  endspecify

endmodule // CMPR42X2TH
`endcelldefine
//$Id: cmpr.genpp,v 1.8 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CMPR42X4TH (S, CO, ICO, A, B, C, D, ICI);
output S, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or  I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor I7 (S, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or  I11 (CO, t5, t6, t7);
  specify
    // delay parameters
    specparam
      tplh$A$S = 1.0,
      tphl$A$S = 1.0,
      tplh$B$S = 1.0,
      tphl$B$S = 1.0,
      tplh$C$S = 1.0,
      tphl$C$S = 1.0,
      tplh$D$S = 1.0,
      tphl$D$S = 1.0,
      tplh$ICI$S = 1.0,
      tphl$ICI$S = 1.0,
      tplh$A$CO = 1.0,
      tphl$A$CO = 1.0,
      tplh$B$CO = 1.0,
      tphl$B$CO = 1.0,
      tplh$C$CO = 1.0,
      tphl$C$CO = 1.0,
      tplh$D$CO = 1.0,
      tphl$D$CO = 1.0,
      tplh$ICI$CO = 1.0,
      tphl$ICI$CO = 1.0,
      tplh$A$ICO = 1.0,
      tphl$A$ICO = 1.0,
      tplh$B$ICO = 1.0,
      tphl$B$ICO = 1.0,
      tplh$C$ICO = 1.0,
      tphl$C$ICO = 1.0,
      tplh$D$ICO = 1.0,
      tphl$D$ICO = 1.0,
      tplh$ICI$ICO = 1.0,
      tphl$ICI$ICO = 1.0;
    // path delays
     if (B == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) 
	(A *> S) = (tplh$A$S, tphl$A$S);
     if (!(B == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) )
	(A *> S) = (tplh$A$S, tphl$A$S);
     if (A == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) 
	(B *> S) = (tplh$B$S, tphl$B$S);
     if (!(A == 1'b1 ^ C == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1) )
	(B *> S) = (tplh$B$S, tphl$B$S);
     if (A == 1'b1 ^ B == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1)
	(C *> S) = (tplh$C$S, tphl$C$S);
     if (!(A == 1'b1 ^ B == 1'b1 ^ D == 1'b1 ^ ICI == 1'b1))
	(C *> S) = (tplh$C$S, tphl$C$S);
     if (A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ ICI == 1'b1)
	(D *> S) = (tplh$D$S, tphl$D$S);
     if (!(A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ ICI == 1'b1))
	(D *> S) = (tplh$D$S, tphl$D$S);
     if (A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ D == 1'b1)
	(ICI *> S) = (tplh$ICI$S, tphl$ICI$S);
     if (!(A == 1'b1 ^ B == 1'b1 ^ C == 1'b1 ^ D == 1'b1))
	(ICI *> S) = (tplh$ICI$S, tphl$ICI$S);
    if (B == 1'b1 && C == 1'b0 )
       (A *> ICO) = (tplh$A$ICO, tphl$A$ICO); 
    if (B == 1'b0 && C == 1'b1 )
       (A *> ICO) = (tplh$A$ICO, tphl$A$ICO); 
    if (A == 1'b1 && C == 1'b0 )
       (B *> ICO) = (tplh$B$ICO, tphl$B$ICO); 
    if (A == 1'b0 && C == 1'b1 )
       (B *> ICO) = (tplh$B$ICO, tphl$B$ICO); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> ICO) = (tplh$C$ICO, tphl$C$ICO); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> ICO) = (tplh$C$ICO, tphl$C$ICO); 
    if (B == 1'b0 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b1 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b0 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && C == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && C == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && C == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && B == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b1 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b0 && D == 1'b1 && ICI == 1'b0 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b1 && B == 1'b0 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b1 && D == 1'b0 && ICI == 1'b1 )
       (C *> CO) = (tplh$C$CO, tphl$C$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && ICI == 1'b1 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && ICI == 1'b0 )
       (D *> CO) = (tplh$D$CO, tphl$D$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO); 
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0 )
       (ICI *> CO) = (tplh$ICI$CO, tphl$ICI$CO);
 
  endspecify

endmodule // CMPR42X4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFX1TH ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFX1TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFX2TH ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFX4TH ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFXLTH ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFXLTH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFHX1TH ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFHX1TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFHX2TH ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFHX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFHX4TH ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFHX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFHXLTH ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFHXLTH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDHX1TH ( S, CO, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0;


     if (B == 1'b1)
	(A *> S) = (tplh$A$S,  tphl$A$S);
     if (B == 1'b0)
	(A *> S)  = (tplh$A$S,  tphl$A$S);
     if (A == 1'b1)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     if (A == 1'b0)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     (A *> CO) = (tplh$A$CO, tphl$A$CO);
     (B *> CO) = (tplh$B$CO, tphl$B$CO);

  endspecify
endmodule // ADDHX1TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDHX2TH ( S, CO, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0;


     if (B == 1'b1)
	(A *> S) = (tplh$A$S,  tphl$A$S);
     if (B == 1'b0)
	(A *> S)  = (tplh$A$S,  tphl$A$S);
     if (A == 1'b1)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     if (A == 1'b0)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     (A *> CO) = (tplh$A$CO, tphl$A$CO);
     (B *> CO) = (tplh$B$CO, tphl$B$CO);

  endspecify
endmodule // ADDHX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDHX4TH ( S, CO, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0;


     if (B == 1'b1)
	(A *> S) = (tplh$A$S,  tphl$A$S);
     if (B == 1'b0)
	(A *> S)  = (tplh$A$S,  tphl$A$S);
     if (A == 1'b1)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     if (A == 1'b0)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     (A *> CO) = (tplh$A$CO, tphl$A$CO);
     (B *> CO) = (tplh$B$CO, tphl$B$CO);

  endspecify
endmodule // ADDHX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDHXLTH ( S, CO, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0;


     if (B == 1'b1)
	(A *> S) = (tplh$A$S,  tphl$A$S);
     if (B == 1'b0)
	(A *> S)  = (tplh$A$S,  tphl$A$S);
     if (A == 1'b1)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     if (A == 1'b0)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     (A *> CO) = (tplh$A$CO, tphl$A$CO);
     (B *> CO) = (tplh$B$CO, tphl$B$CO);

  endspecify
endmodule // ADDHXLTH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AFCSHCINX2TH ( S, CO0, CO1, A, B, CI0N, CI1N, CS);
output S, CO0, CO1;
input A, B, CI0N, CI1N, CS;
  not I0 (cin1, CI1N);
  not I1 (cin0, CI0N);
  xor I2 (s1, A, B, cin1);
  xor I3 (s2, A, B, cin0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or  I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, cin0);
  and I10 (b_and_ci0, B, cin0);
  or  I11 (CO0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, cin1);
  and I13 (b_and_ci1, B, cin1);
  or  I14 (CO1, a_and_b, a_and_ci1, b_and_ci1);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO0  = 1.0,
      tphl$A$CO0  = 1.0,
      tplh$A$CO1  = 1.0,
      tphl$A$CO1  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO0  = 1.0,
      tphl$B$CO0  = 1.0,
      tplh$B$CO1  = 1.0,
      tphl$B$CO1  = 1.0,
      tplh$CI0N$S  = 1.0,
      tphl$CI0N$S  = 1.0,
      tplh$CI0N$CO0  = 1.0,
      tphl$CI0N$CO0  = 1.0,
      tplh$CI0N$CO1  = 1.0,
      tphl$CI0N$CO1  = 1.0,
      tplh$CI1N$S  = 1.0,
      tphl$CI1N$S  = 1.0,
      tplh$CI1N$CO0  = 1.0,
      tphl$CI1N$CO0  = 1.0,
      tplh$CI1N$CO1  = 1.0,
      tphl$CI1N$CO1  = 1.0,
      tplh$CS$S  = 1.0,
      tphl$CS$S  = 1.0,
      tplh$CS$CO0  = 1.0,
      tphl$CS$CO0  = 1.0,
      tplh$CS$CO1  = 1.0,
      tphl$CS$CO1  = 1.0;


    if (A == 1'b1 && B == 1'b0 )
       (CI1N *> CO1) = (tplh$CI1N$CO1, tphl$CI1N$CO1); 
    if (A == 1'b0 && B == 1'b1 )
       (CI1N *> CO1) = (tplh$CI1N$CO1, tphl$CI1N$CO1); 
    if (A == 1'b1 && CI1N == 1'b1 )
       (B *> CO1) = (tplh$B$CO1, tphl$B$CO1); 
    if (A == 1'b0 && CI1N == 1'b0 )
       (B *> CO1) = (tplh$B$CO1, tphl$B$CO1); 
    if (B == 1'b1 && CI1N == 1'b1 )
       (A *> CO1) = (tplh$A$CO1, tphl$A$CO1); 
    if (B == 1'b0 && CI1N == 1'b0 )
       (A *> CO1) = (tplh$A$CO1, tphl$A$CO1); 
    if (A == 1'b1 && CI0N == 1'b1 )
       (B *> CO0) = (tplh$B$CO0, tphl$B$CO0); 
    if (A == 1'b0 && CI0N == 1'b0 )
       (B *> CO0) = (tplh$B$CO0, tphl$B$CO0); 
    if (B == 1'b1 && CI0N == 1'b1 )
       (A *> CO0) = (tplh$A$CO0, tphl$A$CO0); 
    if (B == 1'b0 && CI0N == 1'b0 )
       (A *> CO0) = (tplh$A$CO0, tphl$A$CO0); 
    if (A == 1'b1 && B == 1'b0 )
       (CI0N *> CO0) = (tplh$CI0N$CO0, tphl$CI0N$CO0); 
    if (A == 1'b0 && B == 1'b1 )
       (CI0N *> CO0) = (tplh$CI0N$CO0, tphl$CI0N$CO0); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b0 && CI0N == 1'b1 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b1 && CI0N == 1'b1 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b0 && CI0N == 1'b0 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b1 && CI0N == 1'b0 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b1 && CI0N == 1'b1 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b0 && CI0N == 1'b1 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b1 && CI0N == 1'b0 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b0 && CI0N == 1'b0 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1N == 1'b1 && CI0N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1N == 1'b0 && CI0N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1N == 1'b0 && CI0N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1N == 1'b0 && CI0N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1N == 1'b0 && CI0N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0N == 1'b1 && CI1N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0N == 1'b1 && CI1N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1N == 1'b1 && CI0N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0N == 1'b1 && CI1N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0N == 1'b1 && CI1N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0N == 1'b0 && CI1N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0N == 1'b0 && CI1N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1N == 1'b1 && CI0N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1N == 1'b1 && CI0N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0N == 1'b0 && CI1N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0N == 1'b0 && CI1N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1N == 1'b1 && CI0N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1N == 1'b1 && CI0N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1N == 1'b1 && CI0N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1N == 1'b1 && CI0N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0N == 1'b0 && CI1N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0N == 1'b0 && CI1N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1N == 1'b0 && CI0N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1N == 1'b0 && CI0N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0N == 1'b1 && CI1N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0N == 1'b0 && CI1N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0N == 1'b0 && CI1N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0N == 1'b1 && CI1N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1N == 1'b0 && CI0N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1N == 1'b0 && CI0N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0N == 1'b1 && CI1N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0N == 1'b1 && CI1N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b0 && CI1N == 1'b1 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b1 && CI1N == 1'b1 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b1 && CI1N == 1'b1 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b0 && CI1N == 1'b1 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b1 && CI1N == 1'b0 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b0 && CI1N == 1'b0 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b0 && CI1N == 1'b0 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b1 && CI1N == 1'b0 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (A == 1'b0 && B == 1'b0 && CI0N == 1'b1 && CI1N == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b1 && CI0N == 1'b1 && CI1N == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b1 && CI0N == 1'b0 && CI1N == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b0 && CI0N == 1'b1 && CI1N == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b0 && CI0N == 1'b0 && CI1N == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b0 && CI0N == 1'b0 && CI1N == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b1 && CI0N == 1'b0 && CI1N == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b1 && CI0N == 1'b1 && CI1N == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S);

  endspecify
endmodule // AFCSHCINX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AFCSHCINX4TH ( S, CO0, CO1, A, B, CI0N, CI1N, CS);
output S, CO0, CO1;
input A, B, CI0N, CI1N, CS;
  not I0 (cin1, CI1N);
  not I1 (cin0, CI0N);
  xor I2 (s1, A, B, cin1);
  xor I3 (s2, A, B, cin0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or  I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, cin0);
  and I10 (b_and_ci0, B, cin0);
  or  I11 (CO0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, cin1);
  and I13 (b_and_ci1, B, cin1);
  or  I14 (CO1, a_and_b, a_and_ci1, b_and_ci1);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO0  = 1.0,
      tphl$A$CO0  = 1.0,
      tplh$A$CO1  = 1.0,
      tphl$A$CO1  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO0  = 1.0,
      tphl$B$CO0  = 1.0,
      tplh$B$CO1  = 1.0,
      tphl$B$CO1  = 1.0,
      tplh$CI0N$S  = 1.0,
      tphl$CI0N$S  = 1.0,
      tplh$CI0N$CO0  = 1.0,
      tphl$CI0N$CO0  = 1.0,
      tplh$CI0N$CO1  = 1.0,
      tphl$CI0N$CO1  = 1.0,
      tplh$CI1N$S  = 1.0,
      tphl$CI1N$S  = 1.0,
      tplh$CI1N$CO0  = 1.0,
      tphl$CI1N$CO0  = 1.0,
      tplh$CI1N$CO1  = 1.0,
      tphl$CI1N$CO1  = 1.0,
      tplh$CS$S  = 1.0,
      tphl$CS$S  = 1.0,
      tplh$CS$CO0  = 1.0,
      tphl$CS$CO0  = 1.0,
      tplh$CS$CO1  = 1.0,
      tphl$CS$CO1  = 1.0;


    if (A == 1'b1 && B == 1'b0 )
       (CI1N *> CO1) = (tplh$CI1N$CO1, tphl$CI1N$CO1); 
    if (A == 1'b0 && B == 1'b1 )
       (CI1N *> CO1) = (tplh$CI1N$CO1, tphl$CI1N$CO1); 
    if (A == 1'b1 && CI1N == 1'b1 )
       (B *> CO1) = (tplh$B$CO1, tphl$B$CO1); 
    if (A == 1'b0 && CI1N == 1'b0 )
       (B *> CO1) = (tplh$B$CO1, tphl$B$CO1); 
    if (B == 1'b1 && CI1N == 1'b1 )
       (A *> CO1) = (tplh$A$CO1, tphl$A$CO1); 
    if (B == 1'b0 && CI1N == 1'b0 )
       (A *> CO1) = (tplh$A$CO1, tphl$A$CO1); 
    if (A == 1'b1 && CI0N == 1'b1 )
       (B *> CO0) = (tplh$B$CO0, tphl$B$CO0); 
    if (A == 1'b0 && CI0N == 1'b0 )
       (B *> CO0) = (tplh$B$CO0, tphl$B$CO0); 
    if (B == 1'b1 && CI0N == 1'b1 )
       (A *> CO0) = (tplh$A$CO0, tphl$A$CO0); 
    if (B == 1'b0 && CI0N == 1'b0 )
       (A *> CO0) = (tplh$A$CO0, tphl$A$CO0); 
    if (A == 1'b1 && B == 1'b0 )
       (CI0N *> CO0) = (tplh$CI0N$CO0, tphl$CI0N$CO0); 
    if (A == 1'b0 && B == 1'b1 )
       (CI0N *> CO0) = (tplh$CI0N$CO0, tphl$CI0N$CO0); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b0 && CI0N == 1'b1 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b1 && CI0N == 1'b1 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b0 && CI0N == 1'b0 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b1 && CI0N == 1'b0 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b1 && CI0N == 1'b1 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b0 && CI0N == 1'b1 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b1 && CI0N == 1'b0 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b0 && CI0N == 1'b0 )
       (CI1N *> S) = (tplh$CI1N$S, tphl$CI1N$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1N == 1'b1 && CI0N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1N == 1'b0 && CI0N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1N == 1'b0 && CI0N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1N == 1'b0 && CI0N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1N == 1'b0 && CI0N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0N == 1'b1 && CI1N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0N == 1'b1 && CI1N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1N == 1'b1 && CI0N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0N == 1'b1 && CI1N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0N == 1'b1 && CI1N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0N == 1'b0 && CI1N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0N == 1'b0 && CI1N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1N == 1'b1 && CI0N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1N == 1'b1 && CI0N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0N == 1'b0 && CI1N == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0N == 1'b0 && CI1N == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1N == 1'b1 && CI0N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1N == 1'b1 && CI0N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1N == 1'b1 && CI0N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1N == 1'b1 && CI0N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0N == 1'b0 && CI1N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0N == 1'b0 && CI1N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1N == 1'b0 && CI0N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1N == 1'b0 && CI0N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0N == 1'b1 && CI1N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0N == 1'b0 && CI1N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0N == 1'b0 && CI1N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0N == 1'b1 && CI1N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1N == 1'b0 && CI0N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1N == 1'b0 && CI0N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0N == 1'b1 && CI1N == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0N == 1'b1 && CI1N == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b0 && CI1N == 1'b1 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b1 && CI1N == 1'b1 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b1 && CI1N == 1'b1 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b0 && CI1N == 1'b1 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b1 && CI1N == 1'b0 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b0 && CI1N == 1'b0 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b0 && CI1N == 1'b0 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b1 && CI1N == 1'b0 )
       (CI0N *> S) = (tplh$CI0N$S, tphl$CI0N$S); 
    if (A == 1'b0 && B == 1'b0 && CI0N == 1'b1 && CI1N == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b1 && CI0N == 1'b1 && CI1N == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b1 && CI0N == 1'b0 && CI1N == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b0 && CI0N == 1'b1 && CI1N == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b0 && CI0N == 1'b0 && CI1N == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b0 && CI0N == 1'b0 && CI1N == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b1 && CI0N == 1'b0 && CI1N == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b1 && CI0N == 1'b1 && CI1N == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S);

  endspecify
endmodule // AFCSHCINX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AFCSHCONX2TH ( S, CO0N, CO1N, A, B, CI0, CI1, CS);
output S, CO0N, CO1N;
input A, B, CI0, CI1, CS;
  xor I2 (s1, A, B, CI1);
  xor I3 (s2, A, B, CI0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or  I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, CI0);
  and I10 (b_and_ci0, B, CI0);
  or  I11 (cout0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, CI1);
  and I13 (b_and_ci1, B, CI1);
  or  I14 (cout1, a_and_b, a_and_ci1, b_and_ci1);
  not I15 (CO0N, cout0);
  not I16 (CO1N, cout1);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO0N  = 1.0,
      tphl$A$CO0N  = 1.0,
      tplh$A$CO1N  = 1.0,
      tphl$A$CO1N  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO0N  = 1.0,
      tphl$B$CO0N  = 1.0,
      tplh$B$CO1N  = 1.0,
      tphl$B$CO1N  = 1.0,
      tplh$CI0$S  = 1.0,
      tphl$CI0$S  = 1.0,
      tplh$CI0$CO0N  = 1.0,
      tphl$CI0$CO0N  = 1.0,
      tplh$CI0$CO1N  = 1.0,
      tphl$CI0$CO1N  = 1.0,
      tplh$CI1$S  = 1.0,
      tphl$CI1$S  = 1.0,
      tplh$CI1$CO0N  = 1.0,
      tphl$CI1$CO0N  = 1.0,
      tplh$CI1$CO1N  = 1.0,
      tphl$CI1$CO1N  = 1.0,
      tplh$CS$S  = 1.0,
      tphl$CS$S  = 1.0,
      tplh$CS$CO0N  = 1.0,
      tphl$CS$CO0N  = 1.0,
      tplh$CS$CO1N  = 1.0,
      tphl$CS$CO1N  = 1.0;


    if (CS == 1'b1 && A == 1'b0 && CI1 == 1'b0 && CI0 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1 == 1'b0 && CI0 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1 == 1'b0 && CI0 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1 == 1'b0 && CI0 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1 == 1'b1 && CI0 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1 == 1'b1 && CI0 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1 == 1'b1 && CI0 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1 == 1'b1 && CI0 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CI0 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CI0 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CI0 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CI0 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CI0 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CI0 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CI0 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CI0 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b0 && CI1 == 1'b0 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b1 && CI1 == 1'b0 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b0 && CI1 == 1'b0 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b1 && CI1 == 1'b1 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b0 && CI1 == 1'b1 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b1 && CI1 == 1'b0 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b0 && CI1 == 1'b1 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b1 && CI1 == 1'b1 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b0 && CI0 == 1'b0 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b1 && CI0 == 1'b1 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b1 && CI0 == 1'b0 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b0 && CI0 == 1'b0 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b1 && CI0 == 1'b1 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b0 && CI0 == 1'b1 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b1 && CI0 == 1'b0 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b0 && CI0 == 1'b1 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && CI0 == 1'b0 )
       (B *> CO0N) = (tplh$B$CO0N, tphl$B$CO0N); 
    if (A == 1'b0 && CI0 == 1'b1 )
       (B *> CO0N) = (tplh$B$CO0N, tphl$B$CO0N); 
    if (B == 1'b1 && CI0 == 1'b0 )
       (A *> CO0N) = (tplh$A$CO0N, tphl$A$CO0N); 
    if (B == 1'b0 && CI0 == 1'b1 )
       (A *> CO0N) = (tplh$A$CO0N, tphl$A$CO0N); 
    if (A == 1'b1 && B == 1'b0 )
       (CI0 *> CO0N) = (tplh$CI0$CO0N, tphl$CI0$CO0N); 
    if (A == 1'b0 && B == 1'b1 )
       (CI0 *> CO0N) = (tplh$CI0$CO0N, tphl$CI0$CO0N); 
    if (A == 1'b1 && CI1 == 1'b0 )
       (B *> CO1N) = (tplh$B$CO1N, tphl$B$CO1N); 
    if (A == 1'b0 && CI1 == 1'b1 )
       (B *> CO1N) = (tplh$B$CO1N, tphl$B$CO1N); 
    if (B == 1'b1 && CI1 == 1'b0 )
       (A *> CO1N) = (tplh$A$CO1N, tphl$A$CO1N); 
    if (B == 1'b0 && CI1 == 1'b1 )
       (A *> CO1N) = (tplh$A$CO1N, tphl$A$CO1N); 
    if (A == 1'b1 && B == 1'b0 )
       (CI1 *> CO1N) = (tplh$CI1$CO1N, tphl$CI1$CO1N); 
    if (A == 1'b0 && B == 1'b1 )
       (CI1 *> CO1N) = (tplh$CI1$CO1N, tphl$CI1$CO1N);

  endspecify
endmodule // AFCSHCONX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AFCSHCONX4TH ( S, CO0N, CO1N, A, B, CI0, CI1, CS);
output S, CO0N, CO1N;
input A, B, CI0, CI1, CS;
  xor I2 (s1, A, B, CI1);
  xor I3 (s2, A, B, CI0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or  I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, CI0);
  and I10 (b_and_ci0, B, CI0);
  or  I11 (cout0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, CI1);
  and I13 (b_and_ci1, B, CI1);
  or  I14 (cout1, a_and_b, a_and_ci1, b_and_ci1);
  not I15 (CO0N, cout0);
  not I16 (CO1N, cout1);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO0N  = 1.0,
      tphl$A$CO0N  = 1.0,
      tplh$A$CO1N  = 1.0,
      tphl$A$CO1N  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO0N  = 1.0,
      tphl$B$CO0N  = 1.0,
      tplh$B$CO1N  = 1.0,
      tphl$B$CO1N  = 1.0,
      tplh$CI0$S  = 1.0,
      tphl$CI0$S  = 1.0,
      tplh$CI0$CO0N  = 1.0,
      tphl$CI0$CO0N  = 1.0,
      tplh$CI0$CO1N  = 1.0,
      tphl$CI0$CO1N  = 1.0,
      tplh$CI1$S  = 1.0,
      tphl$CI1$S  = 1.0,
      tplh$CI1$CO0N  = 1.0,
      tphl$CI1$CO0N  = 1.0,
      tplh$CI1$CO1N  = 1.0,
      tphl$CI1$CO1N  = 1.0,
      tplh$CS$S  = 1.0,
      tphl$CS$S  = 1.0,
      tplh$CS$CO0N  = 1.0,
      tphl$CS$CO0N  = 1.0,
      tplh$CS$CO1N  = 1.0,
      tphl$CS$CO1N  = 1.0;


    if (CS == 1'b1 && A == 1'b0 && CI1 == 1'b0 && CI0 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1 == 1'b0 && CI0 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1 == 1'b0 && CI0 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1 == 1'b0 && CI0 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1 == 1'b1 && CI0 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b1 && CI1 == 1'b1 && CI0 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1 == 1'b1 && CI0 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && A == 1'b0 && CI1 == 1'b1 && CI0 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b0 && A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 )
       (B *> S) = (tplh$B$S, tphl$B$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CI0 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CI0 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CI0 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CI0 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CI0 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CI0 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CI0 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CI0 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b0 && CI1 == 1'b0 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b1 && CI1 == 1'b0 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b0 && CI1 == 1'b0 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b1 && CI1 == 1'b1 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b0 && CI1 == 1'b1 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b1 && CI1 == 1'b0 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b0 && B == 1'b0 && CI1 == 1'b1 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b0 && A == 1'b1 && B == 1'b1 && CI1 == 1'b1 )
       (CI0 *> S) = (tplh$CI0$S, tphl$CI0$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b0 && CI0 == 1'b0 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b1 && CI0 == 1'b1 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b1 && CI0 == 1'b0 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b0 && CI0 == 1'b0 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b1 && CI0 == 1'b1 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b0 && CI0 == 1'b1 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b1 && B == 1'b1 && CI0 == 1'b0 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (CS == 1'b1 && A == 1'b0 && B == 1'b0 && CI0 == 1'b1 )
       (CI1 *> S) = (tplh$CI1$S, tphl$CI1$S); 
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && CI0 == 1'b0 )
       (B *> CO0N) = (tplh$B$CO0N, tphl$B$CO0N); 
    if (A == 1'b0 && CI0 == 1'b1 )
       (B *> CO0N) = (tplh$B$CO0N, tphl$B$CO0N); 
    if (B == 1'b1 && CI0 == 1'b0 )
       (A *> CO0N) = (tplh$A$CO0N, tphl$A$CO0N); 
    if (B == 1'b0 && CI0 == 1'b1 )
       (A *> CO0N) = (tplh$A$CO0N, tphl$A$CO0N); 
    if (A == 1'b1 && B == 1'b0 )
       (CI0 *> CO0N) = (tplh$CI0$CO0N, tphl$CI0$CO0N); 
    if (A == 1'b0 && B == 1'b1 )
       (CI0 *> CO0N) = (tplh$CI0$CO0N, tphl$CI0$CO0N); 
    if (A == 1'b1 && CI1 == 1'b0 )
       (B *> CO1N) = (tplh$B$CO1N, tphl$B$CO1N); 
    if (A == 1'b0 && CI1 == 1'b1 )
       (B *> CO1N) = (tplh$B$CO1N, tphl$B$CO1N); 
    if (B == 1'b1 && CI1 == 1'b0 )
       (A *> CO1N) = (tplh$A$CO1N, tphl$A$CO1N); 
    if (B == 1'b0 && CI1 == 1'b1 )
       (A *> CO1N) = (tplh$A$CO1N, tphl$A$CO1N); 
    if (A == 1'b1 && B == 1'b0 )
       (CI1 *> CO1N) = (tplh$CI1$CO1N, tphl$CI1$CO1N); 
    if (A == 1'b0 && B == 1'b1 )
       (CI1 *> CO1N) = (tplh$CI1$CO1N, tphl$CI1$CO1N);

  endspecify
endmodule // AFCSHCONX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AFCSIHCONX2TH ( S, CO0N, CO1N, A, B, CS);
output S, CO0N, CO1N;
input A, B, CS;
  xor I0 (S, A, B, CS);
  and I1 (CO0, A, B);
  or  I2 (CO1, A, B);
  not I3 (CO0N, CO0);
  not I4 (CO1N, CO1);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO0N  = 1.0,
      tphl$A$CO0N  = 1.0,
      tplh$A$CO1N  = 1.0,
      tphl$A$CO1N  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO0N  = 1.0,
      tphl$B$CO0N  = 1.0,
      tplh$B$CO1N  = 1.0,
      tphl$B$CO1N  = 1.0,
      tplh$CS$S  = 1.0,
      tphl$CS$S  = 1.0,
      tplh$CS$CO0N  = 1.0,
      tphl$CS$CO0N  = 1.0,
      tplh$CS$CO1N  = 1.0,
      tphl$CS$CO1N  = 1.0;


     if (B == 1'b0 && CS == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CS == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CS == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CS == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CS == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CS == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
	(A  *> CO0N)  = (tplh$A$CO0N,   tphl$A$CO0N);
	(B  *> CO0N)  = (tplh$B$CO0N,   tphl$B$CO0N);
	(A  *> CO1N)  = (tplh$A$CO1N,   tphl$A$CO1N);
	(B  *> CO1N)  = (tplh$B$CO1N,   tphl$B$CO1N);
    if (A == 1'b0 && B == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S);

  endspecify
endmodule // AFCSIHCONX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AFCSIHCONX4TH ( S, CO0N, CO1N, A, B, CS);
output S, CO0N, CO1N;
input A, B, CS;
  xor I0 (S, A, B, CS);
  and I1 (CO0, A, B);
  or  I2 (CO1, A, B);
  not I3 (CO0N, CO0);
  not I4 (CO1N, CO1);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO0N  = 1.0,
      tphl$A$CO0N  = 1.0,
      tplh$A$CO1N  = 1.0,
      tphl$A$CO1N  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO0N  = 1.0,
      tphl$B$CO0N  = 1.0,
      tplh$B$CO1N  = 1.0,
      tphl$B$CO1N  = 1.0,
      tplh$CS$S  = 1.0,
      tphl$CS$S  = 1.0,
      tplh$CS$CO0N  = 1.0,
      tphl$CS$CO0N  = 1.0,
      tplh$CS$CO1N  = 1.0,
      tphl$CS$CO1N  = 1.0;


     if (B == 1'b0 && CS == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CS == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CS == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CS == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CS == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CS == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
	(A  *> CO0N)  = (tplh$A$CO0N,   tphl$A$CO0N);
	(B  *> CO0N)  = (tplh$B$CO0N,   tphl$B$CO0N);
	(A  *> CO1N)  = (tplh$A$CO1N,   tphl$A$CO1N);
	(B  *> CO1N)  = (tplh$B$CO1N,   tphl$B$CO1N);
    if (A == 1'b0 && B == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CS *> S) = (tplh$CS$S, tphl$CS$S);

  endspecify
endmodule // AFCSIHCONX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AFHCINX2TH ( S, CO, A, B, CIN);
output S, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (S, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or  I5 (CO, a_and_b, a_and_ci, b_and_ci);   
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CIN$S  = 1.0,
      tphl$CIN$S  = 1.0,
      tplh$CIN$CO  = 1.0,
      tphl$CIN$CO  = 1.0;


     if (B == 1'b0 && CIN == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CIN == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CIN == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CIN == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CIN == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CIN == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CIN == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CIN == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
    if (A == 1'b0 && B == 1'b0 )
       (CIN *> S) = (tplh$CIN$S, tphl$CIN$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CIN *> S) = (tplh$CIN$S, tphl$CIN$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CIN *> S) = (tplh$CIN$S, tphl$CIN$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CIN *> S) = (tplh$CIN$S, tphl$CIN$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CIN *> CO) = (tplh$CIN$CO, tphl$CIN$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CIN *> CO) = (tplh$CIN$CO, tphl$CIN$CO); 
    if (A == 1'b1 && CIN == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CIN == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (B == 1'b1 && CIN == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CIN == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO);

  endspecify
endmodule // AFHCINX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AFHCINX4TH ( S, CO, A, B, CIN);
output S, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (S, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or  I5 (CO, a_and_b, a_and_ci, b_and_ci);   
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CIN$S  = 1.0,
      tphl$CIN$S  = 1.0,
      tplh$CIN$CO  = 1.0,
      tphl$CIN$CO  = 1.0;


     if (B == 1'b0 && CIN == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CIN == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CIN == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CIN == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CIN == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CIN == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CIN == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CIN == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
    if (A == 1'b0 && B == 1'b0 )
       (CIN *> S) = (tplh$CIN$S, tphl$CIN$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CIN *> S) = (tplh$CIN$S, tphl$CIN$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CIN *> S) = (tplh$CIN$S, tphl$CIN$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CIN *> S) = (tplh$CIN$S, tphl$CIN$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CIN *> CO) = (tplh$CIN$CO, tphl$CIN$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CIN *> CO) = (tplh$CIN$CO, tphl$CIN$CO); 
    if (A == 1'b1 && CIN == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CIN == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (B == 1'b1 && CIN == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CIN == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO);

  endspecify
endmodule // AFHCINX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AFHCONX2TH ( S, CON, A, B, CI);
output S, CON;
input A, B, CI;
  xor I0 (S, A, B, CI);
  and I1 (a_and_b, A, B);
  and I2 (a_and_ci, A, CI);
  and I3 (b_and_ci, B, CI);
  or  I4 (cout, a_and_b, a_and_ci, b_and_ci);   
  not I5 (CON, cout);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CON  = 1.0,
      tphl$A$CON  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CON  = 1.0,
      tphl$B$CON  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CON  = 1.0,
      tphl$CI$CON  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CON) = (tplh$A$CON, tphl$A$CON); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CON) = (tplh$A$CON, tphl$A$CON); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CON) = (tplh$B$CON, tphl$B$CON); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CON) = (tplh$B$CON, tphl$B$CON); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CON) = (tplh$CI$CON, tphl$CI$CON); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CON) = (tplh$CI$CON, tphl$CI$CON); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // AFHCONX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AFHCONX4TH ( S, CON, A, B, CI);
output S, CON;
input A, B, CI;
  xor I0 (S, A, B, CI);
  and I1 (a_and_b, A, B);
  and I2 (a_and_ci, A, CI);
  and I3 (b_and_ci, B, CI);
  or  I4 (cout, a_and_b, a_and_ci, b_and_ci);   
  not I5 (CON, cout);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CON  = 1.0,
      tphl$A$CON  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CON  = 1.0,
      tphl$B$CON  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CON  = 1.0,
      tphl$CI$CON  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CON) = (tplh$A$CON, tphl$A$CON); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CON) = (tplh$A$CON, tphl$A$CON); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CON) = (tplh$B$CON, tphl$B$CON); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CON) = (tplh$B$CON, tphl$B$CON); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CON) = (tplh$CI$CON, tphl$CI$CON); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CON) = (tplh$CI$CON, tphl$CI$CON); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // AFHCONX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AHCSHCINX2TH ( S, CO, A, CIN, CS);
output S, CO;
input A, CIN, CS;
  not I0 (ci, CIN);
  not I1 (csn, CS);
  xor I2 (s1, A, ci);
  and I3 (s2, CS, s1);
  and I4 (s3, A, csn);
  or  I5 (S, s2, s3);
  and I6 (CO, A, ci);   
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$CIN$S  = 1.0,
      tphl$CIN$S  = 1.0,
      tplh$CIN$CO  = 1.0,
      tphl$CIN$CO  = 1.0,
      tplh$CS$S  = 1.0,
      tphl$CS$S  = 1.0,
      tplh$CS$CO  = 1.0,
      tphl$CS$CO  = 1.0;


     if (A == 1'b0 && CIN == 1'b0)
	(CS  *> S)  = (tplh$CS$S,   tphl$CS$S);
     if (A == 1'b1 && CIN == 1'b0)
	(CS  *> S)  = (tplh$CS$S,   tphl$CS$S);
     if (CIN == 1'b0 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (CIN == 1'b1 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b1 && CS == 1'b1) 
	(CIN  *> S)  = (tplh$CIN$S,   tphl$CIN$S);
     if (A == 1'b0 && CS == 1'b1) 
	(CIN  *> S)  = (tplh$CIN$S,   tphl$CIN$S);
     (A  *> CO)  = (tplh$A$CO,   tphl$A$CO);
     (CIN  *> CO)  = (tplh$CIN$CO,   tphl$CIN$CO);
    if (CIN == 1'b0 && CS == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CIN == 1'b1 && CS == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S);

  endspecify
endmodule // AHCSHCINX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AHCSHCINX4TH ( S, CO, A, CIN, CS);
output S, CO;
input A, CIN, CS;
  not I0 (ci, CIN);
  not I1 (csn, CS);
  xor I2 (s1, A, ci);
  and I3 (s2, CS, s1);
  and I4 (s3, A, csn);
  or  I5 (S, s2, s3);
  and I6 (CO, A, ci);   
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$CIN$S  = 1.0,
      tphl$CIN$S  = 1.0,
      tplh$CIN$CO  = 1.0,
      tphl$CIN$CO  = 1.0,
      tplh$CS$S  = 1.0,
      tphl$CS$S  = 1.0,
      tplh$CS$CO  = 1.0,
      tphl$CS$CO  = 1.0;


     if (A == 1'b0 && CIN == 1'b0)
	(CS  *> S)  = (tplh$CS$S,   tphl$CS$S);
     if (A == 1'b1 && CIN == 1'b0)
	(CS  *> S)  = (tplh$CS$S,   tphl$CS$S);
     if (CIN == 1'b0 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (CIN == 1'b1 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b1 && CS == 1'b1) 
	(CIN  *> S)  = (tplh$CIN$S,   tphl$CIN$S);
     if (A == 1'b0 && CS == 1'b1) 
	(CIN  *> S)  = (tplh$CIN$S,   tphl$CIN$S);
     (A  *> CO)  = (tplh$A$CO,   tphl$A$CO);
     (CIN  *> CO)  = (tplh$CIN$CO,   tphl$CIN$CO);
    if (CIN == 1'b0 && CS == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CIN == 1'b1 && CS == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S);

  endspecify
endmodule // AHCSHCINX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AHCSHCONX2TH ( S, CON, A, CI, CS);
output S, CON;
input A, CI, CS;
  not I1 (csn, CS);
  xor I2 (s1, A, CI);
  and I3 (s2, CS, s1);
  and I4 (s3, A, csn);
  or I5 (S, s2, s3);
  and I6 (cout, A, CI);   
  not I0 (CON, cout);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CON  = 1.0,
      tphl$A$CON  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CON  = 1.0,
      tphl$CI$CON  = 1.0,
      tplh$CS$S  = 1.0,
      tphl$CS$S  = 1.0,
      tplh$CS$CON  = 1.0,
      tphl$CS$CON  = 1.0;


     if (A == 1'b0 && CI == 1'b1)
	(CS  *> S)  = (tplh$CS$S,   tphl$CS$S);
     if (A == 1'b1 && CI == 1'b1)
	(CS  *> S)  = (tplh$CS$S,   tphl$CS$S);
     if (CI == 1'b0 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (CI == 1'b1 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b1 && CS == 1'b1) 
	(CI  *> S)  = (tplh$CI$S,   tphl$CI$S);
     if (A == 1'b0 && CS == 1'b1) 
	(CI  *> S)  = (tplh$CI$S,   tphl$CI$S);
     (A  *> CON)  = (tplh$A$CON,   tphl$A$CON);
     (CI  *> CON)  = (tplh$CI$CON,   tphl$CI$CON);

    if (CI == 1'b1 && CS == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CI == 1'b0 && CS == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S);

  endspecify
endmodule // AHCSHCONX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AHCSHCONX4TH ( S, CON, A, CI, CS);
output S, CON;
input A, CI, CS;
  not I1 (csn, CS);
  xor I2 (s1, A, CI);
  and I3 (s2, CS, s1);
  and I4 (s3, A, csn);
  or I5 (S, s2, s3);
  and I6 (cout, A, CI);   
  not I0 (CON, cout);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CON  = 1.0,
      tphl$A$CON  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CON  = 1.0,
      tphl$CI$CON  = 1.0,
      tplh$CS$S  = 1.0,
      tphl$CS$S  = 1.0,
      tplh$CS$CON  = 1.0,
      tphl$CS$CON  = 1.0;


     if (A == 1'b0 && CI == 1'b1)
	(CS  *> S)  = (tplh$CS$S,   tphl$CS$S);
     if (A == 1'b1 && CI == 1'b1)
	(CS  *> S)  = (tplh$CS$S,   tphl$CS$S);
     if (CI == 1'b0 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (CI == 1'b1 && CS == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b1 && CS == 1'b1) 
	(CI  *> S)  = (tplh$CI$S,   tphl$CI$S);
     if (A == 1'b0 && CS == 1'b1) 
	(CI  *> S)  = (tplh$CI$S,   tphl$CI$S);
     (A  *> CON)  = (tplh$A$CON,   tphl$A$CON);
     (CI  *> CON)  = (tplh$CI$CON,   tphl$CI$CON);

    if (CI == 1'b1 && CS == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S); 
    if (CI == 1'b0 && CS == 1'b0 )
       (A *> S) = (tplh$A$S, tphl$A$S);

  endspecify
endmodule // AHCSHCONX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AHHCINX2TH ( S, CO, A, CIN);
output S, CO;
input A, CIN;
  not I0 (ci, CIN);
  xor I1 (S, A, ci);
  and I2 (CO, A, ci);   
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$CIN$S  = 1.0,
      tphl$CIN$S  = 1.0,
      tplh$CIN$CO  = 1.0,
      tphl$CIN$CO  = 1.0;


    if (CIN == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
    if (CIN == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
    if (A == 1'b1)
	(CIN  *> S)  = (tplh$CIN$S,   tphl$CIN$S);
    if (A == 1'b0)
	(CIN  *> S)  = (tplh$CIN$S,   tphl$CIN$S);
    (A  *> CO)  = (tplh$A$CO,   tphl$A$CO);
    (CIN *> CO) = (tplh$CIN$CO, tphl$CIN$CO);

  endspecify
endmodule // AHHCINX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AHHCINX4TH ( S, CO, A, CIN);
output S, CO;
input A, CIN;
  not I0 (ci, CIN);
  xor I1 (S, A, ci);
  and I2 (CO, A, ci);   
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$CIN$S  = 1.0,
      tphl$CIN$S  = 1.0,
      tplh$CIN$CO  = 1.0,
      tphl$CIN$CO  = 1.0;


    if (CIN == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
    if (CIN == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
    if (A == 1'b1)
	(CIN  *> S)  = (tplh$CIN$S,   tphl$CIN$S);
    if (A == 1'b0)
	(CIN  *> S)  = (tplh$CIN$S,   tphl$CIN$S);
    (A  *> CO)  = (tplh$A$CO,   tphl$A$CO);
    (CIN *> CO) = (tplh$CIN$CO, tphl$CIN$CO);

  endspecify
endmodule // AHHCINX4TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AHHCONX2TH ( S, CON, A, CI);
output S, CON;
input A, CI;
  xor I0 (S, A, CI);
  and  I1 (cout, A, CI);   
  not I2 (CON, cout);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CON  = 1.0,
      tphl$A$CON  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CON  = 1.0,
      tphl$CI$CON  = 1.0;


    if (CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
    if (CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
    if (A == 1'b1)
	(CI  *> S)  = (tplh$CI$S,   tphl$CI$S);
    if (A == 1'b0)
	(CI  *> S)  = (tplh$CI$S,   tphl$CI$S);
    (A  *> CON)  = (tplh$A$CON,   tphl$A$CON);
    (CI *> CON) = (tplh$CI$CON, tphl$CI$CON);

  endspecify
endmodule // AHHCONX2TH
`endcelldefine
//$Id: add.genpp,v 1.6 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AHHCONX4TH ( S, CON, A, CI);
output S, CON;
input A, CI;
  xor I0 (S, A, CI);
  and  I1 (cout, A, CI);   
  not I2 (CON, cout);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CON  = 1.0,
      tphl$A$CON  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CON  = 1.0,
      tphl$CI$CON  = 1.0;


    if (CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
    if (CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
    if (A == 1'b1)
	(CI  *> S)  = (tplh$CI$S,   tphl$CI$S);
    if (A == 1'b0)
	(CI  *> S)  = (tplh$CI$S,   tphl$CI$S);
    (A  *> CON)  = (tplh$A$CON,   tphl$A$CON);
    (CI *> CON) = (tplh$CI$CON, tphl$CI$CON);

  endspecify
endmodule // AHHCONX4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X1TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X2TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X4TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X6TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X8TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2XLTH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X1TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X2TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X4TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X6TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X8TH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3XLTH (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X1TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X2TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X4TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X6TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X8TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4XLTH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4XLTH
`endcelldefine
//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X1TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X2TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X4TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21XLTH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X1TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X2TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X4TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22XLTH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO2B2X1TH (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // AO2B2X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO2B2X2TH (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // AO2B2X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO2B2X4TH (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // AO2B2X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO2B2XLTH (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  and I2 (outB, B0, B1);
  or I3 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // AO2B2XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO2B2BX1TH (Y, A0, A1N, B0, B1N);
output Y;
input A0, A1N, B0, B1N;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1N$Y = 1.0,
      tphl$B1N$Y = 1.0;

    // path delays
    if (A1N == 1'b0 && B0 == 1'b1 && B1N == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1N == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1N == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1N == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1N == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (B1N == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1N == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1N == 1'b0 && A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y);

  endspecify
endmodule // AO2B2BX1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO2B2BX2TH (Y, A0, A1N, B0, B1N);
output Y;
input A0, A1N, B0, B1N;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1N$Y = 1.0,
      tphl$B1N$Y = 1.0;

    // path delays
    if (A1N == 1'b0 && B0 == 1'b1 && B1N == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1N == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1N == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1N == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1N == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (B1N == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1N == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1N == 1'b0 && A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y);

  endspecify
endmodule // AO2B2BX2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO2B2BX4TH (Y, A0, A1N, B0, B1N);
output Y;
input A0, A1N, B0, B1N;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1N$Y = 1.0,
      tphl$B1N$Y = 1.0;

    // path delays
    if (A1N == 1'b0 && B0 == 1'b1 && B1N == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1N == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1N == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1N == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1N == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (B1N == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1N == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1N == 1'b0 && A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y);

  endspecify
endmodule // AO2B2BX4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO2B2BXLTH (Y, A0, A1N, B0, B1N);
output Y;
input A0, A1N, B0, B1N;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  not I2 (outB1, B1N);
  and I3 (outB, B0, outB1);
  or I4 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1N$Y = 1.0,
      tphl$B1N$Y = 1.0;

    // path delays
    if (A1N == 1'b0 && B0 == 1'b1 && B1N == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1N == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1N == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1N == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1N == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (B1N == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1N == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1N == 1'b0 && A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1N == 1'b1 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b0 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1N == 1'b1 )
       (B1N *> Y) = (tplh$B1N$Y, tphl$B1N$Y);

  endspecify
endmodule // AO2B2BXLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211X1TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211X2TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211X4TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211XLTH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X1TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X2TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X3TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X3TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X4TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X6TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X6TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X8TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X8TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21XLTH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX1TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX2TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX4TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BXLTH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BXLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221X1TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221X2TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221X4TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221XLTH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222X1TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222X2TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222X4TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222XLTH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X1TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X2TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X4TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22XLTH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2B1X1TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2B1X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2B1X2TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2B1X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2B1X4TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2B1X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2B1XLTH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2B1XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2BB1X1TH (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;

  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2BB1X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2BB1X2TH (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;

  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2BB1X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2BB1X4TH (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;

  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2BB1X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2BB1XLTH (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;

  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2BB1XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2BB2X1TH (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;

  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b1 && A0N == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0N == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0N == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0N == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A0N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // AOI2BB2X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2BB2X2TH (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;

  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b1 && A0N == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0N == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0N == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0N == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A0N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // AOI2BB2X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2BB2X4TH (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;

  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b1 && A0N == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0N == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0N == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0N == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A0N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // AOI2BB2X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2BB2XLTH (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;

  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b1 && A0N == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0N == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0N == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0N == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A0N == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // AOI2BB2XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X1TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X2TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X4TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31XLTH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X1TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X2TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X4TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32XLTH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI33X1TH (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$B2$Y = 1.0,
      tphl$B2$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y);

  endspecify
endmodule // AOI33X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI33X2TH (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$B2$Y = 1.0,
      tphl$B2$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y);

  endspecify
endmodule // AOI33X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI33X4TH (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$B2$Y = 1.0,
      tphl$B2$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y);

  endspecify
endmodule // AOI33X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI33XLTH (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$B2$Y = 1.0,
      tphl$B2$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && B2 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b1 && B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y);

  endspecify
endmodule // AOI33XLTH
`endcelldefine





//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX10TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX10TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX12TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX12TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX14TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX14TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX16TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX16TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX18TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX18TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX20TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX20TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX2TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX2TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX3TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX3TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX4TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX4TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX5TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX5TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX6TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX6TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX8TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKAND2X12TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // CLKAND2X12TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKAND2X2TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // CLKAND2X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKAND2X3TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // CLKAND2X3TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKAND2X4TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // CLKAND2X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKAND2X6TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // CLKAND2X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKAND2X8TH (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // CLKAND2X8TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX12TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX12TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX16TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX16TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX1TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX1TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX20TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX20TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX24TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX24TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX2TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX2TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX32TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX32TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX3TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX3TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX40TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX40TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX4TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX4TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX6TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX6TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKBUFX8TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKBUFX8TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX12TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX12TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX16TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX16TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX1TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX1TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX20TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX20TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX24TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX24TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX2TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX2TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX32TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX32TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX3TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX3TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX40TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX40TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX4TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX4TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX6TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX6TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKINVX8TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // CLKINVX8TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKMX2X12TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKMX2X12TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKMX2X2TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKMX2X2TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKMX2X3TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKMX2X3TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKMX2X4TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKMX2X4TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKMX2X6TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKMX2X6TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKMX2X8TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKMX2X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKNAND2X12TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // CLKNAND2X12TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKNAND2X2TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // CLKNAND2X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKNAND2X4TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // CLKNAND2X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKNAND2X8TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // CLKNAND2X8TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKXOR2X12TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKXOR2X12TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKXOR2X1TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKXOR2X1TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKXOR2X2TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKXOR2X2TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKXOR2X4TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKXOR2X4TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module CLKXOR2X8TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // CLKXOR2X8TH
`endcelldefine
//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFX1TH (Q, QN, D, CK);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFX2TH (Q, QN, D, CK);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFX4TH (Q, QN, D, CK);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFXLTH (Q, QN, D, CK);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFXLTH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFHX1TH (Q, QN, D, CK);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFHX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFHX2TH (Q, QN, D, CK);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFHX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFHX4TH (Q, QN, D, CK);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFHX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFHX8TH (Q, QN, D, CK);
output Q, QN;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFHX8TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFHQX1TH (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFHQX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFHQX2TH (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFHQX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFHQX4TH (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFHQX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFHQX8TH (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFHQX8TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNHX1TH (Q, QN, D, CKN);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tplh$CKN$QN	= 1.0,
    tphl$CKN$QN	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (flag)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);

   endspecify
endmodule // DFFNHX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNHX2TH (Q, QN, D, CKN);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tplh$CKN$QN	= 1.0,
    tphl$CKN$QN	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (flag)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);

   endspecify
endmodule // DFFNHX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNHX4TH (Q, QN, D, CKN);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tplh$CKN$QN	= 1.0,
    tphl$CKN$QN	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (flag)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);

   endspecify
endmodule // DFFNHX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNHX8TH (Q, QN, D, CKN);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
wire dD;
wire dCKN;
supply1 xSN,xRN;
supply1 dSN, dRN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tplh$CKN$QN	= 1.0,
    tphl$CKN$QN	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (flag)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);

   endspecify
endmodule // DFFNHX8TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNSRHX1TH (Q, QN, D, CKN, SN, RN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tplh$CKN$QN	= 1.0,
    tphl$CKN$QN	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tsetup$SN$CKN    = 1.0,
    thold$SN$CKN    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CKN    = 1.0,
    thold$RN$CKN    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (flag)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN, posedge RN &&& (SN == 1'b1), tsetup$RN$CKN, thold$RN$CKN, NOTIFIER, , ,dCKN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN, thold$SN$CKN, NOTIFIER, , ,dCKN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFNSRHX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNSRHX2TH (Q, QN, D, CKN, SN, RN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tplh$CKN$QN	= 1.0,
    tphl$CKN$QN	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tsetup$SN$CKN    = 1.0,
    thold$SN$CKN    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CKN    = 1.0,
    thold$RN$CKN    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (flag)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN, posedge RN &&& (SN == 1'b1), tsetup$RN$CKN, thold$RN$CKN, NOTIFIER, , ,dCKN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN, thold$SN$CKN, NOTIFIER, , ,dCKN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFNSRHX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNSRHX4TH (Q, QN, D, CKN, SN, RN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tplh$CKN$QN	= 1.0,
    tphl$CKN$QN	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tsetup$SN$CKN    = 1.0,
    thold$SN$CKN    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CKN    = 1.0,
    thold$RN$CKN    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (flag)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN, posedge RN &&& (SN == 1'b1), tsetup$RN$CKN, thold$RN$CKN, NOTIFIER, , ,dCKN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN, thold$SN$CKN, NOTIFIER, , ,dCKN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFNSRHX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNSRHX8TH (Q, QN, D, CKN, SN, RN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tplh$CKN$QN	= 1.0,
    tphl$CKN$QN	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tsetup$SN$CKN    = 1.0,
    thold$SN$CKN    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CKN    = 1.0,
    thold$RN$CKN    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (flag)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN, posedge RN &&& (SN == 1'b1), tsetup$RN$CKN, thold$RN$CKN, NOTIFIER, , ,dCKN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN, thold$SN$CKN, NOTIFIER, , ,dCKN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFNSRHX8TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQX1TH (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQX2TH (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQX4TH (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQXLTH (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQXLTH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRX1TH (Q, QN, D, CK, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFRX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRX2TH (Q, QN, D, CK, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFRX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRX4TH (Q, QN, D, CK, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFRX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRXLTH (Q, QN, D, CK, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFRXLTH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRHQX1TH (Q, D, CK, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFRHQX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRHQX2TH (Q, D, CK, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFRHQX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRHQX4TH (Q, D, CK, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFRHQX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRHQX8TH (Q, D, CK, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFRHQX8TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRQX1TH (Q, D, CK, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFRQX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRQX2TH (Q, D, CK, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFRQX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRQX4TH (Q, D, CK, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFRQX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRQXLTH (Q, D, CK, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN;

  buf   XX0 (xRN, RN);
supply1 dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFRQXLTH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSX1TH (Q, QN, D, CK, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule // DFFSX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSX2TH (Q, QN, D, CK, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule // DFFSX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSX4TH (Q, QN, D, CK, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule // DFFSX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSXLTH (Q, QN, D, CK, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule // DFFSXLTH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSHQX1TH (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSHQX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSHQX2TH (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSHQX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSHQX4TH (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSHQX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSHQX8TH (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSHQX8TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQX1TH (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSQX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQX2TH (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSQX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQX4TH (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSQX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQXLTH (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
supply1 xRN;

  buf   XX0 (xSN, SN);
supply1 dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSQXLTH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRX1TH (Q, QN, D, CK, SN, RN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFSRX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRX2TH (Q, QN, D, CK, SN, RN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFSRX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRX4TH (Q, QN, D, CK, SN, RN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFSRX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRXLTH (Q, QN, D, CK, SN, RN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

   endspecify
endmodule // DFFSRXLTH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRHQX1TH (Q, D, CK, SN, RN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFSRHQX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRHQX2TH (Q, D, CK, SN, RN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFSRHQX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRHQX4TH (Q, D, CK, SN, RN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFSRHQX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRHQX8TH (Q, D, CK, SN, RN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$RN$CK    = 1.0,
    thold$RN$CK    = 0.5,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    thold$RN$SN = 1.0,
    thold$SN$RN = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK, thold$RN$CK, NOTIFIER, , , dCK, dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER, , , dCK, dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && RN == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule // DFFSRHQX8TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFTRX1TH (Q, QN, D, CK, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
supply1 dSN, dEN;
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, dCK);
  udp_edfft I0 (n0, dD, clk, dRN, dSN, dEN, NOTIFIER);
  buf     I1 (Q, n0);
  and     I4 (Deff, dD, dRN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$RN$CK = 0.5,
    tsetup$RN$CK = 1.0,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    (posedge CK *> (Q  +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
    (posedge CK *> (QN -: Deff)) = (tplh$CK$QN, tphl$CK$QN);
 
    // timing checks
    $setuphold(posedge CK &&& (rn_and_sn == 1), posedge D,  tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (rn_and_sn == 1), negedge D,  tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (xSN == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $setuphold(posedge CK &&& (xSN == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFTRX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFTRX2TH (Q, QN, D, CK, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
supply1 dSN, dEN;
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, dCK);
  udp_edfft I0 (n0, dD, clk, dRN, dSN, dEN, NOTIFIER);
  buf     I1 (Q, n0);
  and     I4 (Deff, dD, dRN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$RN$CK = 0.5,
    tsetup$RN$CK = 1.0,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    (posedge CK *> (Q  +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
    (posedge CK *> (QN -: Deff)) = (tplh$CK$QN, tphl$CK$QN);
 
    // timing checks
    $setuphold(posedge CK &&& (rn_and_sn == 1), posedge D,  tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (rn_and_sn == 1), negedge D,  tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (xSN == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $setuphold(posedge CK &&& (xSN == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFTRX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFTRX4TH (Q, QN, D, CK, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
supply1 dSN, dEN;
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, dCK);
  udp_edfft I0 (n0, dD, clk, dRN, dSN, dEN, NOTIFIER);
  buf     I1 (Q, n0);
  and     I4 (Deff, dD, dRN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$RN$CK = 0.5,
    tsetup$RN$CK = 1.0,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    (posedge CK *> (Q  +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
    (posedge CK *> (QN -: Deff)) = (tplh$CK$QN, tphl$CK$QN);
 
    // timing checks
    $setuphold(posedge CK &&& (rn_and_sn == 1), posedge D,  tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (rn_and_sn == 1), negedge D,  tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (xSN == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $setuphold(posedge CK &&& (xSN == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFTRX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFTRXLTH (Q, QN, D, CK, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dRN;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
supply1 dSN, dEN;
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, dCK);
  udp_edfft I0 (n0, dD, clk, dRN, dSN, dEN, NOTIFIER);
  buf     I1 (Q, n0);
  and     I4 (Deff, dD, dRN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$RN$Q  = 1.0,
    tphl$RN$Q  = 1.0,
    tplh$RN$QN  = 1.0,
    tphl$RN$QN  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$RN$CK = 0.5,
    tsetup$RN$CK = 1.0,
    tminpwl$RN     = 1.0,
    tminpwh$RN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    (posedge CK *> (Q  +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
    (posedge CK *> (QN -: Deff)) = (tplh$CK$QN, tphl$CK$QN);
 
    // timing checks
    $setuphold(posedge CK &&& (rn_and_sn == 1), posedge D,  tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (rn_and_sn == 1), negedge D,  tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (xSN == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $setuphold(posedge CK &&& (xSN == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFTRXLTH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFYQX2TH (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
wire dD;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
  and     I4 (flag, dRN, dSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFYQX2TH
`endcelldefine


//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DLY1X1TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // DLY1X1TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DLY1X4TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // DLY1X4TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DLY2X1TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // DLY2X1TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DLY2X4TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // DLY2X4TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DLY3X1TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // DLY3X1TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DLY3X4TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // DLY3X4TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DLY4X1TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // DLY4X1TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DLY4X4TH (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // DLY4X4TH
`endcelldefine
//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFX1TH (Q, QN, D, CK, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);
  and      I2 (flag, dRN, dSN);
  and      I3 (Dcheck, dSN, dRN, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
        (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFX1TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFX2TH (Q, QN, D, CK, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);
  and      I2 (flag, dRN, dSN);
  and      I3 (Dcheck, dSN, dRN, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
        (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFX2TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFX4TH (Q, QN, D, CK, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);
  and      I2 (flag, dRN, dSN);
  and      I3 (Dcheck, dSN, dRN, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
        (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFX4TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFXLTH (Q, QN, D, CK, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);
  and      I2 (flag, dRN, dSN);
  and      I3 (Dcheck, dSN, dRN, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
        (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFXLTH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFHQX1TH (Q, D, CK, E);
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  and      I2 (flag, dRN, dSN);
  and      I3 (Dcheck, dSN, dRN, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFHQX1TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFHQX2TH (Q, D, CK, E);
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  and      I2 (flag, dRN, dSN);
  and      I3 (Dcheck, dSN, dRN, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFHQX2TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFHQX4TH (Q, D, CK, E);
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  and      I2 (flag, dRN, dSN);
  and      I3 (Dcheck, dSN, dRN, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFHQX4TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFHQX8TH (Q, D, CK, E);
output Q;
input D, CK, E;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, dD, dCK, dRN, dSN, dE, NOTIFIER);
  buf     B1 (Q, n0);
  and      I2 (flag, dRN, dSN);
  and      I3 (Dcheck, dSN, dRN, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFHQX8TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFTRX1TH (Q, QN, D, CK, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, dD, dCK, dRN, dSN, E, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  and     I3 (Deff, dRN, dD);
  and     I4 (Dcheck,dE,dRN);
  and     I5 (check,dE, dD);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
    (posedge CK *> (Q  +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
    (posedge CK *> (QN -: Deff)) = (tplh$CK$QN, tphl$CK$QN);   
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge E &&& (RN == 1), tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E &&& (RN == 1), tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $setuphold(posedge CK, negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFTRX1TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFTRX2TH (Q, QN, D, CK, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, dD, dCK, dRN, dSN, E, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  and     I3 (Deff, dRN, dD);
  and     I4 (Dcheck,dE,dRN);
  and     I5 (check,dE, dD);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
    (posedge CK *> (Q  +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
    (posedge CK *> (QN -: Deff)) = (tplh$CK$QN, tphl$CK$QN);   
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge E &&& (RN == 1), tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E &&& (RN == 1), tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $setuphold(posedge CK, negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFTRX2TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFTRX4TH (Q, QN, D, CK, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, dD, dCK, dRN, dSN, E, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  and     I3 (Deff, dRN, dD);
  and     I4 (Dcheck,dE,dRN);
  and     I5 (check,dE, dD);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
    (posedge CK *> (Q  +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
    (posedge CK *> (QN -: Deff)) = (tplh$CK$QN, tphl$CK$QN);   
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge E &&& (RN == 1), tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E &&& (RN == 1), tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $setuphold(posedge CK, negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFTRX4TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFTRXLTH (Q, QN, D, CK, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, dD, dCK, dRN, dSN, E, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);
  and     I3 (Deff, dRN, dD);
  and     I4 (Dcheck,dE,dRN);
  and     I5 (check,dE, dD);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
    (posedge CK *> (Q  +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
    (posedge CK *> (QN -: Deff)) = (tplh$CK$QN, tphl$CK$QN);   
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK, posedge E &&& (RN == 1), tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E &&& (RN == 1), tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
    $setuphold(posedge CK, negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFTRXLTH
`endcelldefine


//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX10TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX10TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX12TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX12TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX14TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX14TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX16TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX16TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX18TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX18TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX1TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX1TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX20TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX20TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX2TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX2TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX3TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX3TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX4TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX4TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX5TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX5TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX6TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX6TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX8TH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX8TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVXLTH (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVXLTH
`endcelldefine
//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MDFFHQX1TH (Q, D0, D1, S0, CK);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff  I1 (n0, nm, clk, dRN, dSN, NOTIFIER);
  not      I2 (nsel,dS0);
  and      I3 (flag0, dRN, dSN, nsel);
  and      I4 (flag1, dRN, dSN, dS0);
  buf      I5 (Q, n0);
  xor      I6 (D0xorD1, dD0, dD1);
  and      I7 (flag, D0xorD1, dRN, dSN);
  and      I8 (SandR,dRN, dSN);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (Q +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag1)
      (posedge CK *> (Q +: D1)) = (tplh$CK$Q,    tphl$CK$Q);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER, , ,dCK,dS0);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER, , ,dCK,dS0);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // MDFFHQX1TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MDFFHQX2TH (Q, D0, D1, S0, CK);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff  I1 (n0, nm, clk, dRN, dSN, NOTIFIER);
  not      I2 (nsel,dS0);
  and      I3 (flag0, dRN, dSN, nsel);
  and      I4 (flag1, dRN, dSN, dS0);
  buf      I5 (Q, n0);
  xor      I6 (D0xorD1, dD0, dD1);
  and      I7 (flag, D0xorD1, dRN, dSN);
  and      I8 (SandR,dRN, dSN);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (Q +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag1)
      (posedge CK *> (Q +: D1)) = (tplh$CK$Q,    tphl$CK$Q);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER, , ,dCK,dS0);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER, , ,dCK,dS0);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // MDFFHQX2TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MDFFHQX4TH (Q, D0, D1, S0, CK);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff  I1 (n0, nm, clk, dRN, dSN, NOTIFIER);
  not      I2 (nsel,dS0);
  and      I3 (flag0, dRN, dSN, nsel);
  and      I4 (flag1, dRN, dSN, dS0);
  buf      I5 (Q, n0);
  xor      I6 (D0xorD1, dD0, dD1);
  and      I7 (flag, D0xorD1, dRN, dSN);
  and      I8 (SandR,dRN, dSN);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (Q +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag1)
      (posedge CK *> (Q +: D1)) = (tplh$CK$Q,    tphl$CK$Q);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER, , ,dCK,dS0);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER, , ,dCK,dS0);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // MDFFHQX4TH
`endcelldefine


//$Id: dff.genpp,v 1.13 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MDFFHQX8TH (Q, D0, D1, S0, CK);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dCK;
supply1 xSN,xRN;
supply1 dSN, dRN;
  buf     IC (clk, dCK);
  udp_mux2 I0 (nm, dD0, dD1, dS0);
  udp_dff  I1 (n0, nm, clk, dRN, dSN, NOTIFIER);
  not      I2 (nsel,dS0);
  and      I3 (flag0, dRN, dSN, nsel);
  and      I4 (flag1, dRN, dSN, dS0);
  buf      I5 (Q, n0);
  xor      I6 (D0xorD1, dD0, dD1);
  and      I7 (flag, D0xorD1, dRN, dSN);
  and      I8 (SandR,dRN, dSN);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (Q +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag1)
      (posedge CK *> (Q +: D1)) = (tplh$CK$Q,    tphl$CK$Q);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER, , ,dCK,dS0);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER, , ,dCK,dS0);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // MDFFHQX8TH
`endcelldefine


//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X1TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X1TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X2TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X2TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X3TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X3TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X4TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X4TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X6TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X6TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X8TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X8TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2XLTH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2XLTH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX3X1TH (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(Y, A, B, C, C, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MX3X1TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX3X2TH (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(Y, A, B, C, C, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MX3X2TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX3X4TH (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(Y, A, B, C, C, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MX3X4TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX3XLTH (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(Y, A, B, C, C, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MX3XLTH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX4X1TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MX4X1TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX4X2TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MX4X2TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX4X4TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MX4X4TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX4XLTH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MX4XLTH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2X1TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2X1TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2X2TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2X2TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2X3TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2X3TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2X4TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2X4TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2X6TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2X6TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2X8TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2X8TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2XLTH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2XLTH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2DX1TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2DX1TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2DX2TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2DX2TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2DX4TH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2DX4TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI2DXLTH (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXI2DXLTH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI3X1TH (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXI3X1TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI3X2TH (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXI3X2TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI3X4TH (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXI3X4TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI3XLTH (Y, A, B, C, S0, S1);
output Y;
input A, B, C, S0, S1;

  udp_mux4 u0(YN,A, B, C, C, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b0 && S0 == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b0 && B == 1'b0 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b1 && S0 == 1'b1 && B == 1'b1 && A == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXI3XLTH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI4X1TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXI4X1TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI4X2TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXI4X2TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI4X4TH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXI4X4TH
`endcelldefine
//$Id: mux.genpp,v 1.8 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXI4XLTH (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXI4XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X1TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X2TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X3TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X3TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X4TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X5TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X5TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X6TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X8TH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2XLTH (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX1TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX2TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX4TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX8TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BXLTH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BXLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X1TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X2TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X3TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X3TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X4TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X6TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X8TH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3XLTH (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX1TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX2TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX4TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BXLTH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BXLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X1TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X2TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X4TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X6TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X8TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4XLTH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BX1TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BX1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BX2TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BX2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BX4TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BX4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BXLTH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BXLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BBX1TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BBX1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BBX2TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BBX2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BBX4TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BBX4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BBXLTH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BBXLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X1TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X2TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X3TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X3TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X4TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X5TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X5TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X6TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X8TH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2XLTH (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX1TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX2TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX4TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX8TH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BXLTH (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BXLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X1TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X2TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X4TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X6TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X8TH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3XLTH (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3BX1TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3BX1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3BX2TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3BX2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3BX4TH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3BX4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3BXLTH (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3BXLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4X1TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4X2TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4X4TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4X6TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4X8TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4XLTH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4BX1TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4BX1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4BX2TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4BX2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4BX4TH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4BX4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4BXLTH (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4BXLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4BBX1TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4BBX1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4BBX2TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4BBX2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4BBX4TH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4BBX4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR4BBXLTH (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NOR4BBXLTH
`endcelldefine
//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X1TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X2TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X4TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21XLTH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X1TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X2TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X4TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22XLTH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211X1TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211X2TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211X4TH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211XLTH (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X1TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X2TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X3TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X3TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X4TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X6TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X6TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X8TH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X8TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21XLTH (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX1TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX2TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX4TH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BXLTH (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BXLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221X1TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221X2TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221X4TH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221XLTH (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222X1TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222X2TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222X4TH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222XLTH (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X1TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X2TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X4TH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22XLTH (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B11X1TH (Y, A0, A1N, B0, C0);
output Y;
input A0, A1N, B0, C0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, outA, B0, C0);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI2B11X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B11X2TH (Y, A0, A1N, B0, C0);
output Y;
input A0, A1N, B0, C0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, outA, B0, C0);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI2B11X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B11X4TH (Y, A0, A1N, B0, C0);
output Y;
input A0, A1N, B0, C0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, outA, B0, C0);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI2B11X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B11XLTH (Y, A0, A1N, B0, C0);
output Y;
input A0, A1N, B0, C0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, outA, B0, C0);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI2B11XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B1X1TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2B1X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B1X2TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2B1X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B1X4TH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2B1X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B1XLTH (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2B1XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B2X1TH (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI2B2X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B2X2TH (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI2B2X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B2X4TH (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI2B2X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2B2XLTH (Y, A0, A1N, B0, B1);
output Y;
input A0, A1N, B0, B1;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  or I2 (outB, B0, B1);
  nand I3 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI2B2XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2BB1X1TH (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;

  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2BB1X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2BB1X2TH (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;

  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2BB1X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2BB1X4TH (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;

  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2BB1X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2BB1XLTH (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;

  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0N == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2BB1XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2BB2X1TH (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;

  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b0 && A0N == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0N == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0N == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0N == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A0N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // OAI2BB2X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2BB2X2TH (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;

  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b0 && A0N == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0N == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0N == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0N == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A0N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // OAI2BB2X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2BB2X4TH (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;

  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b0 && A0N == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0N == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0N == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0N == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A0N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // OAI2BB2X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2BB2XLTH (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;

  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (B1 == 1'b0 && A0N == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0N == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0N == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0N == 1'b0 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0N == 1'b1 && A1N == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0N == 1'b0 && A1N == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A1N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0N *> Y) = (tplh$A0N$Y, tphl$A0N$Y); 
    if (A0N == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y); 
    if (A0N == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);

  endspecify
endmodule // OAI2BB2XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI31X1TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI31X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI31X2TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI31X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI31X4TH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI31X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI31XLTH (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI31XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI32X1TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI32X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI32X2TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI32X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI32X4TH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI32X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI32XLTH (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI32XLTH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI33X1TH (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;

  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$B2$Y = 1.0,
      tphl$B2$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y);

  endspecify
endmodule // OAI33X1TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI33X2TH (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;

  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$B2$Y = 1.0,
      tphl$B2$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y);

  endspecify
endmodule // OAI33X2TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI33X4TH (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;

  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$B2$Y = 1.0,
      tphl$B2$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y);

  endspecify
endmodule // OAI33X4TH
`endcelldefine





//$Id: aoi.genpp,v 1.7 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI33XLTH (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;

  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$B2$Y = 1.0,
      tphl$B2$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A2 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b0 && A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && B2 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y); 
    if (B1 == 1'b0 && B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b1 )
       (B2 *> Y) = (tplh$B2$Y, tphl$B2$Y);

  endspecify
endmodule // OAI33XLTH
`endcelldefine





//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X1TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X2TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X4TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X6TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X8TH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2XLTH (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X1TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X2TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X4TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X6TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X8TH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3XLTH (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3XLTH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X1TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X1TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X2TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X2TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X4TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X4TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X6TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X6TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X8TH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X8TH
`endcelldefine
//$Id: comb.genpp,v 1.4 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4XLTH (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4XLTH
`endcelldefine
//$Id: bmux.genpp,v 1.8 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BMXX2TH (PP, X2, A, S, M1, M0);
output PP;
input X2, A, S, M1, M0;

  udp_bmx I0 (PP, X2, A, S, M1, M0);
  specify
    // delay parameters
    specparam
      tplh$X2$PP = 1.0,
      tphl$X2$PP = 1.0,
      tplh$A$PP = 1.0,
      tphl$A$PP = 1.0,
      tplh$S$PP = 1.0,
      tphl$S$PP = 1.0,
      tplh$M1$PP = 1.0,
      tphl$M1$PP = 1.0,
      tplh$M0$PP = 1.0,
      tphl$M0$PP = 1.0;
    // path delays
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b1 && M1 == 1'b0 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b1 && M1 == 1'b1 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b1 && M0 == 1'b1 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b0 && M1 == 1'b0 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b0 && M1 == 1'b1 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b1 && M0 == 1'b0 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b0 && M0 == 1'b0 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b0 && M0 == 1'b1 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b1 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b0 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b0 && M0 == 1'b1 && A == 1'b0 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b1 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b0 && M0 == 1'b1 && A == 1'b1 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b0 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b0 && A == 1'b0 && M0 == 1'b0 && S == 1'b1 )
       (M1 *> PP) = (tplh$M1$PP, tphl$M1$PP); 
    if (X2 == 1'b0 && A == 1'b1 && M0 == 1'b0 && S == 1'b0 )
       (M1 *> PP) = (tplh$M1$PP, tphl$M1$PP); 
    if (X2 == 1'b0 && A == 1'b0 && M0 == 1'b1 && S == 1'b1 )
       (M1 *> PP) = (tplh$M1$PP, tphl$M1$PP); 
    if (X2 == 1'b0 && A == 1'b1 && M0 == 1'b1 && S == 1'b0 )
       (M1 *> PP) = (tplh$M1$PP, tphl$M1$PP); 
    if (X2 == 1'b1 && A == 1'b0 && M1 == 1'b0 && S == 1'b1 )
       (M0 *> PP) = (tplh$M0$PP, tphl$M0$PP); 
    if (X2 == 1'b1 && A == 1'b1 && M1 == 1'b0 && S == 1'b0 )
       (M0 *> PP) = (tplh$M0$PP, tphl$M0$PP); 
    if (X2 == 1'b1 && A == 1'b0 && M1 == 1'b1 && S == 1'b1 )
       (M0 *> PP) = (tplh$M0$PP, tphl$M0$PP); 
    if (X2 == 1'b1 && A == 1'b1 && M1 == 1'b1 && S == 1'b0 )
       (M0 *> PP) = (tplh$M0$PP, tphl$M0$PP); 
    if (M0 == 1'b1 && A == 1'b1 && M1 == 1'b0 && S == 1'b0 )
       (X2 *> PP) = (tplh$X2$PP, tphl$X2$PP); 
    if (M0 == 1'b0 && S == 1'b1 && M1 == 1'b1 && A == 1'b0 )
       (X2 *> PP) = (tplh$X2$PP, tphl$X2$PP); 
    if (M0 == 1'b1 && A == 1'b0 && M1 == 1'b0 && S == 1'b1 )
       (X2 *> PP) = (tplh$X2$PP, tphl$X2$PP); 
    if (M0 == 1'b0 && S == 1'b0 && M1 == 1'b1 && A == 1'b1 )
       (X2 *> PP) = (tplh$X2$PP, tphl$X2$PP);
  endspecify

endmodule // BMXX2TH
`endcelldefine
//$Id: bmux.genpp,v 1.8 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BMXX4TH (PP, X2, A, S, M1, M0);
output PP;
input X2, A, S, M1, M0;

  udp_bmx I0 (PP, X2, A, S, M1, M0);
  specify
    // delay parameters
    specparam
      tplh$X2$PP = 1.0,
      tphl$X2$PP = 1.0,
      tplh$A$PP = 1.0,
      tphl$A$PP = 1.0,
      tplh$S$PP = 1.0,
      tphl$S$PP = 1.0,
      tplh$M1$PP = 1.0,
      tphl$M1$PP = 1.0,
      tplh$M0$PP = 1.0,
      tphl$M0$PP = 1.0;
    // path delays
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b1 && M1 == 1'b0 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b1 && M1 == 1'b1 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b1 && M0 == 1'b1 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b0 && M1 == 1'b0 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b0 && M1 == 1'b1 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b1 && M0 == 1'b0 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b0 && M0 == 1'b0 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b0 && M0 == 1'b1 )
       (A *> PP) = (tplh$A$PP, tphl$A$PP); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b1 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b0 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b0 && M0 == 1'b1 && A == 1'b0 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b1 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b0 && M0 == 1'b1 && A == 1'b1 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b0 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b0 )
       (S *> PP) = (tplh$S$PP, tphl$S$PP); 
    if (X2 == 1'b0 && A == 1'b0 && M0 == 1'b0 && S == 1'b1 )
       (M1 *> PP) = (tplh$M1$PP, tphl$M1$PP); 
    if (X2 == 1'b0 && A == 1'b1 && M0 == 1'b0 && S == 1'b0 )
       (M1 *> PP) = (tplh$M1$PP, tphl$M1$PP); 
    if (X2 == 1'b0 && A == 1'b0 && M0 == 1'b1 && S == 1'b1 )
       (M1 *> PP) = (tplh$M1$PP, tphl$M1$PP); 
    if (X2 == 1'b0 && A == 1'b1 && M0 == 1'b1 && S == 1'b0 )
       (M1 *> PP) = (tplh$M1$PP, tphl$M1$PP); 
    if (X2 == 1'b1 && A == 1'b0 && M1 == 1'b0 && S == 1'b1 )
       (M0 *> PP) = (tplh$M0$PP, tphl$M0$PP); 
    if (X2 == 1'b1 && A == 1'b1 && M1 == 1'b0 && S == 1'b0 )
       (M0 *> PP) = (tplh$M0$PP, tphl$M0$PP); 
    if (X2 == 1'b1 && A == 1'b0 && M1 == 1'b1 && S == 1'b1 )
       (M0 *> PP) = (tplh$M0$PP, tphl$M0$PP); 
    if (X2 == 1'b1 && A == 1'b1 && M1 == 1'b1 && S == 1'b0 )
       (M0 *> PP) = (tplh$M0$PP, tphl$M0$PP); 
    if (M0 == 1'b1 && A == 1'b1 && M1 == 1'b0 && S == 1'b0 )
       (X2 *> PP) = (tplh$X2$PP, tphl$X2$PP); 
    if (M0 == 1'b0 && S == 1'b1 && M1 == 1'b1 && A == 1'b0 )
       (X2 *> PP) = (tplh$X2$PP, tphl$X2$PP); 
    if (M0 == 1'b1 && A == 1'b0 && M1 == 1'b0 && S == 1'b1 )
       (X2 *> PP) = (tplh$X2$PP, tphl$X2$PP); 
    if (M0 == 1'b0 && S == 1'b0 && M1 == 1'b1 && A == 1'b1 )
       (X2 *> PP) = (tplh$X2$PP, tphl$X2$PP);
  endspecify

endmodule // BMXX4TH
`endcelldefine
//$Id: bmux.genpp,v 1.8 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BMXIX2TH (PPN, X2, A, S, M1, M0);
output PPN;
input X2, A, S, M1, M0;

  udp_bmx I0 (nPP, X2, A, S, M1, M0);
  not  I1 (PPN, nPP);
  specify
    // delay parameters
    specparam
      tplh$X2$PPN = 1.0,
      tphl$X2$PPN = 1.0,
      tplh$A$PPN = 1.0,
      tphl$A$PPN = 1.0,
      tplh$S$PPN = 1.0,
      tphl$S$PPN = 1.0,
      tplh$M1$PPN = 1.0,
      tphl$M1$PPN = 1.0,
      tplh$M0$PPN = 1.0,
      tphl$M0$PPN = 1.0;
    // path delays
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b1 && M1 == 1'b0 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b1 && M1 == 1'b1 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b1 && M0 == 1'b1 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b0 && M1 == 1'b0 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b0 && M1 == 1'b1 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b1 && M0 == 1'b0 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b0 && M0 == 1'b0 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b0 && M0 == 1'b1 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b1 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b0 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b0 && M0 == 1'b1 && A == 1'b0 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b1 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b0 && M0 == 1'b1 && A == 1'b1 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b0 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b0 && A == 1'b0 && M0 == 1'b0 && S == 1'b1 )
       (M1 *> PPN) = (tplh$M1$PPN, tphl$M1$PPN); 
    if (X2 == 1'b0 && A == 1'b1 && M0 == 1'b0 && S == 1'b0 )
       (M1 *> PPN) = (tplh$M1$PPN, tphl$M1$PPN); 
    if (X2 == 1'b0 && A == 1'b0 && M0 == 1'b1 && S == 1'b1 )
       (M1 *> PPN) = (tplh$M1$PPN, tphl$M1$PPN); 
    if (X2 == 1'b0 && A == 1'b1 && M0 == 1'b1 && S == 1'b0 )
       (M1 *> PPN) = (tplh$M1$PPN, tphl$M1$PPN); 
    if (X2 == 1'b1 && A == 1'b0 && M1 == 1'b0 && S == 1'b1 )
       (M0 *> PPN) = (tplh$M0$PPN, tphl$M0$PPN); 
    if (X2 == 1'b1 && A == 1'b1 && M1 == 1'b0 && S == 1'b0 )
       (M0 *> PPN) = (tplh$M0$PPN, tphl$M0$PPN); 
    if (X2 == 1'b1 && A == 1'b0 && M1 == 1'b1 && S == 1'b1 )
       (M0 *> PPN) = (tplh$M0$PPN, tphl$M0$PPN); 
    if (X2 == 1'b1 && A == 1'b1 && M1 == 1'b1 && S == 1'b0 )
       (M0 *> PPN) = (tplh$M0$PPN, tphl$M0$PPN); 
    if (M0 == 1'b1 && A == 1'b1 && M1 == 1'b0 && S == 1'b0 )
       (X2 *> PPN) = (tplh$X2$PPN, tphl$X2$PPN); 
    if (M0 == 1'b0 && S == 1'b1 && M1 == 1'b1 && A == 1'b0 )
       (X2 *> PPN) = (tplh$X2$PPN, tphl$X2$PPN); 
    if (M0 == 1'b1 && A == 1'b0 && M1 == 1'b0 && S == 1'b1 )
       (X2 *> PPN) = (tplh$X2$PPN, tphl$X2$PPN); 
    if (M0 == 1'b0 && S == 1'b0 && M1 == 1'b1 && A == 1'b1 )
       (X2 *> PPN) = (tplh$X2$PPN, tphl$X2$PPN);
  endspecify

endmodule // BMXIX2TH
`endcelldefine
//$Id: bmux.genpp,v 1.8 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BMXIX4TH (PPN, X2, A, S, M1, M0);
output PPN;
input X2, A, S, M1, M0;

  udp_bmx I0 (nPP, X2, A, S, M1, M0);
  not  I1 (PPN, nPP);
  specify
    // delay parameters
    specparam
      tplh$X2$PPN = 1.0,
      tphl$X2$PPN = 1.0,
      tplh$A$PPN = 1.0,
      tphl$A$PPN = 1.0,
      tplh$S$PPN = 1.0,
      tphl$S$PPN = 1.0,
      tplh$M1$PPN = 1.0,
      tphl$M1$PPN = 1.0,
      tplh$M0$PPN = 1.0,
      tphl$M0$PPN = 1.0;
    // path delays
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b1 && M1 == 1'b0 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b1 && M1 == 1'b1 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b1 && M0 == 1'b1 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b0 && M1 == 1'b0 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b1 && M0 == 1'b1 && S == 1'b0 && M1 == 1'b1 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b1 && M0 == 1'b0 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b0 && M0 == 1'b0 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b0 && M1 == 1'b1 && S == 1'b0 && M0 == 1'b1 )
       (A *> PPN) = (tplh$A$PPN, tphl$A$PPN); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b1 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b0 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b0 && M0 == 1'b1 && A == 1'b0 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b1 && M0 == 1'b0 && A == 1'b1 && M1 == 1'b1 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b0 && M0 == 1'b1 && A == 1'b1 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b0 && M0 == 1'b0 && A == 1'b0 && M1 == 1'b0 )
       (S *> PPN) = (tplh$S$PPN, tphl$S$PPN); 
    if (X2 == 1'b0 && A == 1'b0 && M0 == 1'b0 && S == 1'b1 )
       (M1 *> PPN) = (tplh$M1$PPN, tphl$M1$PPN); 
    if (X2 == 1'b0 && A == 1'b1 && M0 == 1'b0 && S == 1'b0 )
       (M1 *> PPN) = (tplh$M1$PPN, tphl$M1$PPN); 
    if (X2 == 1'b0 && A == 1'b0 && M0 == 1'b1 && S == 1'b1 )
       (M1 *> PPN) = (tplh$M1$PPN, tphl$M1$PPN); 
    if (X2 == 1'b0 && A == 1'b1 && M0 == 1'b1 && S == 1'b0 )
       (M1 *> PPN) = (tplh$M1$PPN, tphl$M1$PPN); 
    if (X2 == 1'b1 && A == 1'b0 && M1 == 1'b0 && S == 1'b1 )
       (M0 *> PPN) = (tplh$M0$PPN, tphl$M0$PPN); 
    if (X2 == 1'b1 && A == 1'b1 && M1 == 1'b0 && S == 1'b0 )
       (M0 *> PPN) = (tplh$M0$PPN, tphl$M0$PPN); 
    if (X2 == 1'b1 && A == 1'b0 && M1 == 1'b1 && S == 1'b1 )
       (M0 *> PPN) = (tplh$M0$PPN, tphl$M0$PPN); 
    if (X2 == 1'b1 && A == 1'b1 && M1 == 1'b1 && S == 1'b0 )
       (M0 *> PPN) = (tplh$M0$PPN, tphl$M0$PPN); 
    if (M0 == 1'b1 && A == 1'b1 && M1 == 1'b0 && S == 1'b0 )
       (X2 *> PPN) = (tplh$X2$PPN, tphl$X2$PPN); 
    if (M0 == 1'b0 && S == 1'b1 && M1 == 1'b1 && A == 1'b0 )
       (X2 *> PPN) = (tplh$X2$PPN, tphl$X2$PPN); 
    if (M0 == 1'b1 && A == 1'b0 && M1 == 1'b0 && S == 1'b1 )
       (X2 *> PPN) = (tplh$X2$PPN, tphl$X2$PPN); 
    if (M0 == 1'b0 && S == 1'b0 && M1 == 1'b1 && A == 1'b1 )
       (X2 *> PPN) = (tplh$X2$PPN, tphl$X2$PPN);
  endspecify

endmodule // BMXIX4TH
`endcelldefine
//$Id: bmux.genpp,v 1.8 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BENCX1TH (S, A, X2, M2, M1, M0);
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (S, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (A, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);
  specify
    // delay parameters
    specparam
      tplh$M2$S = 1.0,
      tphl$M2$S = 1.0,
      tplh$M1$S = 1.0,
      tphl$M1$S = 1.0,
      tplh$M0$S = 1.0,
      tphl$M0$S = 1.0,
      tplh$M2$A = 1.0,
      tphl$M2$A = 1.0,
      tplh$M1$A = 1.0,
      tphl$M1$A = 1.0,
      tplh$M0$A = 1.0,
      tphl$M0$A = 1.0,
      tplh$M2$X2 = 1.0,
      tphl$M2$X2 = 1.0,
      tplh$M1$X2 = 1.0,
      tphl$M1$X2 = 1.0,
      tplh$M0$X2 = 1.0,
      tphl$M0$X2 = 1.0;
    // path delays
     if (M0== 1'b1)
	(M1 *> X2) = (tplh$M1$X2, tphl$M1$X2);
     if (M0== 1'b0)
	(M1 *> X2) = (tplh$M1$X2, tphl$M1$X2);
     if (M1== 1'b1)
	(M0 *> X2) = (tplh$M0$X2, tphl$M0$X2);
     if (M1== 1'b0)
	(M0 *> X2) = (tplh$M0$X2, tphl$M0$X2);
     (M0 *> S) = (tplh$M0$S, tphl$M0$S);
     (M1 *> S) = (tplh$M1$S, tphl$M1$S);
     (M0 *> A) = (tplh$M0$A, tphl$M0$A);
     (M1 *> A) = (tplh$M1$A, tphl$M1$A);
    if (M0 == 1'b0 && M1 == 1'b0 )
       (M2 *> S) = (tplh$M2$S, tphl$M2$S); 
    if (M0 == 1'b1 && M1 == 1'b0 )
       (M2 *> S) = (tplh$M2$S, tphl$M2$S); 
    if (M0 == 1'b0 && M1 == 1'b1 )
       (M2 *> S) = (tplh$M2$S, tphl$M2$S); 
    if (M0 == 1'b1 && M1 == 1'b1 )
       (M2 *> A) = (tplh$M2$A, tphl$M2$A); 
    if (M0 == 1'b0 && M1 == 1'b1 )
       (M2 *> A) = (tplh$M2$A, tphl$M2$A); 
    if (M0 == 1'b1 && M1 == 1'b0 )
       (M2 *> A) = (tplh$M2$A, tphl$M2$A);
  endspecify

endmodule // BENCX1TH
`endcelldefine
//$Id: bmux.genpp,v 1.8 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BENCX2TH (S, A, X2, M2, M1, M0);
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (S, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (A, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);
  specify
    // delay parameters
    specparam
      tplh$M2$S = 1.0,
      tphl$M2$S = 1.0,
      tplh$M1$S = 1.0,
      tphl$M1$S = 1.0,
      tplh$M0$S = 1.0,
      tphl$M0$S = 1.0,
      tplh$M2$A = 1.0,
      tphl$M2$A = 1.0,
      tplh$M1$A = 1.0,
      tphl$M1$A = 1.0,
      tplh$M0$A = 1.0,
      tphl$M0$A = 1.0,
      tplh$M2$X2 = 1.0,
      tphl$M2$X2 = 1.0,
      tplh$M1$X2 = 1.0,
      tphl$M1$X2 = 1.0,
      tplh$M0$X2 = 1.0,
      tphl$M0$X2 = 1.0;
    // path delays
     if (M0== 1'b1)
	(M1 *> X2) = (tplh$M1$X2, tphl$M1$X2);
     if (M0== 1'b0)
	(M1 *> X2) = (tplh$M1$X2, tphl$M1$X2);
     if (M1== 1'b1)
	(M0 *> X2) = (tplh$M0$X2, tphl$M0$X2);
     if (M1== 1'b0)
	(M0 *> X2) = (tplh$M0$X2, tphl$M0$X2);
     (M0 *> S) = (tplh$M0$S, tphl$M0$S);
     (M1 *> S) = (tplh$M1$S, tphl$M1$S);
     (M0 *> A) = (tplh$M0$A, tphl$M0$A);
     (M1 *> A) = (tplh$M1$A, tphl$M1$A);
    if (M0 == 1'b0 && M1 == 1'b0 )
       (M2 *> S) = (tplh$M2$S, tphl$M2$S); 
    if (M0 == 1'b1 && M1 == 1'b0 )
       (M2 *> S) = (tplh$M2$S, tphl$M2$S); 
    if (M0 == 1'b0 && M1 == 1'b1 )
       (M2 *> S) = (tplh$M2$S, tphl$M2$S); 
    if (M0 == 1'b1 && M1 == 1'b1 )
       (M2 *> A) = (tplh$M2$A, tphl$M2$A); 
    if (M0 == 1'b0 && M1 == 1'b1 )
       (M2 *> A) = (tplh$M2$A, tphl$M2$A); 
    if (M0 == 1'b1 && M1 == 1'b0 )
       (M2 *> A) = (tplh$M2$A, tphl$M2$A);
  endspecify

endmodule // BENCX2TH
`endcelldefine
//$Id: bmux.genpp,v 1.8 2006/01/09 06:34:37 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BENCX4TH (S, A, X2, M2, M1, M0);
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (S, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (A, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);
  specify
    // delay parameters
    specparam
      tplh$M2$S = 1.0,
      tphl$M2$S = 1.0,
      tplh$M1$S = 1.0,
      tphl$M1$S = 1.0,
      tplh$M0$S = 1.0,
      tphl$M0$S = 1.0,
      tplh$M2$A = 1.0,
      tphl$M2$A = 1.0,
      tplh$M1$A = 1.0,
      tphl$M1$A = 1.0,
      tplh$M0$A = 1.0,
      tphl$M0$A = 1.0,
      tplh$M2$X2 = 1.0,
      tphl$M2$X2 = 1.0,
      tplh$M1$X2 = 1.0,
      tphl$M1$X2 = 1.0,
      tplh$M0$X2 = 1.0,
      tphl$M0$X2 = 1.0;
    // path delays
     if (M0== 1'b1)
	(M1 *> X2) = (tplh$M1$X2, tphl$M1$X2);
     if (M0== 1'b0)
	(M1 *> X2) = (tplh$M1$X2, tphl$M1$X2);
     if (M1== 1'b1)
	(M0 *> X2) = (tplh$M0$X2, tphl$M0$X2);
     if (M1== 1'b0)
	(M0 *> X2) = (tplh$M0$X2, tphl$M0$X2);
     (M0 *> S) = (tplh$M0$S, tphl$M0$S);
     (M1 *> S) = (tplh$M1$S, tphl$M1$S);
     (M0 *> A) = (tplh$M0$A, tphl$M0$A);
     (M1 *> A) = (tplh$M1$A, tphl$M1$A);
    if (M0 == 1'b0 && M1 == 1'b0 )
       (M2 *> S) = (tplh$M2$S, tphl$M2$S); 
    if (M0 == 1'b1 && M1 == 1'b0 )
       (M2 *> S) = (tplh$M2$S, tphl$M2$S); 
    if (M0 == 1'b0 && M1 == 1'b1 )
       (M2 *> S) = (tplh$M2$S, tphl$M2$S); 
    if (M0 == 1'b1 && M1 == 1'b1 )
       (M2 *> A) = (tplh$M2$A, tphl$M2$A); 
    if (M0 == 1'b0 && M1 == 1'b1 )
       (M2 *> A) = (tplh$M2$A, tphl$M2$A); 
    if (M0 == 1'b1 && M1 == 1'b0 )
       (M2 *> A) = (tplh$M2$A, tphl$M2$A);
  endspecify

endmodule // BENCX4TH
`endcelldefine
//$Id: rf.genpp,v 1.10 2006/03/24 11:24:21 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF2R1WX1TH (R1B, R2B, WB, WW, R1W, R2W);
output R1B, R2B;
input WB, WW, R1W, R2W;
reg NOTIFIER;

   not        I0 (WWN, WW);
   not        I1 (R1WN, R1W);
   not        I2 (R2WN, R2W);
   udp_tlatrf I3 (n0, WB, WW, WWN, NOTIFIER);
   notif1     I4 (R1B, n0, n2);
   notif1     I5 (R2B, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, R1W);
   udp_outrf  I7 (n3, n0, R2WN, R2W);

  specify
    // delay parameters
    specparam
      tplh$WB$R1B = 1.0,
      tphl$WB$R1B = 1.0,
      tplh$WW$R1B = 1.0,
      tphl$WW$R1B = 1.0,
      tplh$R1W$R1B = 1.0,
      tphl$R1W$R1B = 1.0,
      tplh$R2W$R1B = 1.0,
      tphl$R2W$R1B = 1.0,
      tplh$WB$R2B = 1.0,
      tphl$WB$R2B = 1.0,
      tplh$WW$R2B = 1.0,
      tphl$WW$R2B = 1.0,
      tplh$R1W$R2B = 1.0,
      tphl$R1W$R2B = 1.0,
      tplh$R2W$R2B = 1.0,
      tphl$R2W$R2B = 1.0,
    tminpwh$WW    = 1.0,
    tperiod$WW    = 1.0,
    tsetup$WW$WB = 1.0,
    thold$WW$WB  = 0.5;

      // path delays
      ( WW *> R1B) = (tplh$WW$R1B, tphl$WW$R1B);
      ( WW *> R2B) = (tplh$WW$R2B, tphl$WW$R2B);
 
      // timing checks
      $width(posedge WW, tminpwh$WW, 0, NOTIFIER);
      $period(posedge WW, tperiod$WW, NOTIFIER);
      $setuphold(negedge WW, posedge WB, tsetup$WW$WB, thold$WW$WB, NOTIFIER);
      $setuphold(negedge WW, negedge WB, tsetup$WW$WB, thold$WW$WB, NOTIFIER);
    if (WW == 1'b1 && R1W == 1'b1 )
       ( WB *> R2B) = (tplh$WB$R2B, tphl$WB$R2B); 
    if (WW == 1'b1 && R1W == 1'b0 )
       ( WB *> R2B) = (tplh$WB$R2B, tphl$WB$R2B); 
    if (R1W == 1'b1 && R2W == 1'b1 )
       (posedge  WW *> (R2B -: WB)) = (tplh$WW$R2B, tphl$WW$R2B); 
    if (R1W == 1'b0 && R2W == 1'b1 )
       (posedge  WW *> (R2B -: WB)) = (tplh$WW$R2B, tphl$WW$R2B); 
    if (WW == 1'b1 && R1W == 1'b1 )
       ( R2W *> R2B) = (tplh$R2W$R2B, tphl$R2W$R2B); 
    if (WB == 1'b1 && WW == 1'b0 && R1W == 1'b1 )
       ( R2W *> R2B) = (tplh$R2W$R2B, tphl$R2W$R2B); 
    if (WW == 1'b1 && R1W == 1'b0 )
       ( R2W *> R2B) = (tplh$R2W$R2B, tphl$R2W$R2B); 
    if (WB == 1'b1 && WW == 1'b0 && R1W == 1'b0 )
       ( R2W *> R2B) = (tplh$R2W$R2B, tphl$R2W$R2B); 
    if (WB == 1'b0 && WW == 1'b0 && R1W == 1'b1 )
       ( R2W *> R2B) = (tplh$R2W$R2B, tphl$R2W$R2B); 
    if (WB == 1'b0 && WW == 1'b0 && R1W == 1'b0 )
       ( R2W *> R2B) = (tplh$R2W$R2B, tphl$R2W$R2B); 
    if (WW == 1'b1 && R2W == 1'b1 )
       ( WB *> R1B) = (tplh$WB$R1B, tphl$WB$R1B); 
    if (WW == 1'b1 && R2W == 1'b0 )
       ( WB *> R1B) = (tplh$WB$R1B, tphl$WB$R1B); 
    if (R1W == 1'b1 && R2W == 1'b1 )
       (posedge  WW *> (R1B -: WB)) = (tplh$WW$R1B, tphl$WW$R1B); 
    if (R1W == 1'b1 && R2W == 1'b0 )
       (posedge  WW *> (R1B -: WB)) = (tplh$WW$R1B, tphl$WW$R1B); 
    if (WW == 1'b1 && R2W == 1'b1 )
       ( R1W *> R1B) = (tplh$R1W$R1B, tphl$R1W$R1B); 
    if (WW == 1'b1 && R2W == 1'b0 )
       ( R1W *> R1B) = (tplh$R1W$R1B, tphl$R1W$R1B); 
    if (WB == 1'b1 && WW == 1'b0 && R2W == 1'b0 )
       ( R1W *> R1B) = (tplh$R1W$R1B, tphl$R1W$R1B); 
    if (WB == 1'b0 && WW == 1'b0 && R2W == 1'b1 )
       ( R1W *> R1B) = (tplh$R1W$R1B, tphl$R1W$R1B); 
    if (WB == 1'b0 && WW == 1'b0 && R2W == 1'b0 )
       ( R1W *> R1B) = (tplh$R1W$R1B, tphl$R1W$R1B); 
    if (WB == 1'b1 && WW == 1'b0 && R2W == 1'b1 )
       ( R1W *> R1B) = (tplh$R1W$R1B, tphl$R1W$R1B);
 

  endspecify

endmodule // RF2R1WX1TH
`endcelldefine
//$Id: rf.genpp,v 1.10 2006/03/24 11:24:21 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF1R1WX1TH (RB, WB, WW, RW, RWN);
output RB;
input WB, WW, RW, RWN;
reg NOTIFIER;

   not II (wwn,WW);
   udp_tlatrf I0 (n0, WB, WW, wwn, NOTIFIER);
   notif1     I1 (RB, n0, n2);
   udp_outrf  I2 (n2, n0, RWN, RW);

  specify
    // delay parameters
    specparam
      tplh$WB$RB = 1.0,
      tphl$WB$RB = 1.0,
      tplh$WW$RB = 1.0,
      tphl$WW$RB = 1.0,
      tplh$RW$RB = 1.0,
      tphl$RW$RB = 1.0,
      tplh$RWN$RB = 1.0,
      tphl$RWN$RB = 1.0,
    tsetup$WW$WB = 1.0,
    thold$WW$WB  = 0.5,
    tminpwh$WW    = 1.0,
    tperiod$WW    = 1.0;

      // path delays
      ( posedge WW *> (RB -:WB )) = (tplh$WW$RB, tphl$WW$RB);
      ( WB *> RB ) = (tplh$WB$RB, tphl$WB$RB);
      ( RW *> RB ) = (tplh$RW$RB, tphl$RW$RB);
      ( RWN *> RB ) = (tplh$RWN$RB, tphl$RWN$RB);
 
      // timing checks
      $width(posedge WW, tminpwh$WW, 0, NOTIFIER);
      $period(posedge WW, tperiod$WW, NOTIFIER);
      $setuphold(negedge WW, posedge WB, tsetup$WW$WB, thold$WW$WB, NOTIFIER);
      $setuphold(negedge WW, negedge WB, tsetup$WW$WB, thold$WW$WB, NOTIFIER);
 

  endspecify

endmodule // RF1R1WX1TH
`endcelldefine
//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFX1TH (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFX2TH (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFX4TH (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFXLTH (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFXLTH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFHX1TH (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFHX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFHX2TH (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFHX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFHX4TH (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFHX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFHX8TH (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFHX8TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFHQX1TH (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFHQX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFHQX2TH (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFHQX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFHQX4TH (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFHQX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFHQX8TH (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFHQX8TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNHX1TH (Q, QN, D, SI, SE, CKN);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tplh$CKN$QN = 1.0,
      tphl$CKN$QN = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSEb)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    if (SandRandSE)
      (negedge CKN *> (QN -: SI)) = (tplh$CKN$QN, tphl$CKN$QN);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);

endspecify
endmodule // SDFFNHX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNHX2TH (Q, QN, D, SI, SE, CKN);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tplh$CKN$QN = 1.0,
      tphl$CKN$QN = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSEb)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    if (SandRandSE)
      (negedge CKN *> (QN -: SI)) = (tplh$CKN$QN, tphl$CKN$QN);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);

endspecify
endmodule // SDFFNHX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNHX4TH (Q, QN, D, SI, SE, CKN);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tplh$CKN$QN = 1.0,
      tphl$CKN$QN = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSEb)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    if (SandRandSE)
      (negedge CKN *> (QN -: SI)) = (tplh$CKN$QN, tphl$CKN$QN);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);

endspecify
endmodule // SDFFNHX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNHX8TH (Q, QN, D, SI, SE, CKN);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tplh$CKN$QN = 1.0,
      tphl$CKN$QN = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSEb)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    if (SandRandSE)
      (negedge CKN *> (QN -: SI)) = (tplh$CKN$QN, tphl$CKN$QN);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);

endspecify
endmodule // SDFFNHX8TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNSRHX1TH (Q, QN, D, SI, SE, CKN, SN, RN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CKN = 1.0,
      thold$SN$CKN = 0.5,
      tsetup$RN$CKN = 1.0,
      thold$RN$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tplh$CKN$QN = 1.0,
      tphl$CKN$QN = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSEb)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    if (SandRandSE)
      (negedge CKN *> (QN -: SI)) = (tplh$CKN$QN, tphl$CKN$QN);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN ,thold$SN$CKN , NOTIFIER, , ,dCKN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge RN &&& (SN == 1'b1), tsetup$RN$CKN ,thold$RN$CKN , NOTIFIER, , ,dCKN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFNSRHX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNSRHX2TH (Q, QN, D, SI, SE, CKN, SN, RN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CKN = 1.0,
      thold$SN$CKN = 0.5,
      tsetup$RN$CKN = 1.0,
      thold$RN$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tplh$CKN$QN = 1.0,
      tphl$CKN$QN = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSEb)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    if (SandRandSE)
      (negedge CKN *> (QN -: SI)) = (tplh$CKN$QN, tphl$CKN$QN);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN ,thold$SN$CKN , NOTIFIER, , ,dCKN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge RN &&& (SN == 1'b1), tsetup$RN$CKN ,thold$RN$CKN , NOTIFIER, , ,dCKN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFNSRHX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNSRHX4TH (Q, QN, D, SI, SE, CKN, SN, RN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CKN = 1.0,
      thold$SN$CKN = 0.5,
      tsetup$RN$CKN = 1.0,
      thold$RN$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tplh$CKN$QN = 1.0,
      tphl$CKN$QN = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSEb)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    if (SandRandSE)
      (negedge CKN *> (QN -: SI)) = (tplh$CKN$QN, tphl$CKN$QN);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN ,thold$SN$CKN , NOTIFIER, , ,dCKN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge RN &&& (SN == 1'b1), tsetup$RN$CKN ,thold$RN$CKN , NOTIFIER, , ,dCKN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFNSRHX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNSRHX8TH (Q, QN, D, SI, SE, CKN, SN, RN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCKN;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, dCKN);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CKN = 1.0,
      thold$SN$CKN = 0.5,
      tsetup$RN$CKN = 1.0,
      thold$RN$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tplh$CKN$QN = 1.0,
      tphl$CKN$QN = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSEb)
      (negedge CKN *> (QN -: D)) = (tplh$CKN$QN, tphl$CKN$QN);
    if (SandRandSE)
      (negedge CKN *> (QN -: SI)) = (tplh$CKN$QN, tphl$CKN$QN);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER, , ,dCKN,dD);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER, , ,dCKN,dSI);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER, , ,dCKN,dSE);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN ,thold$SN$CKN , NOTIFIER, , ,dCKN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge RN &&& (SN == 1'b1), tsetup$RN$CKN ,thold$RN$CKN , NOTIFIER, , ,dCKN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFNSRHX8TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQX1TH (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQX2TH (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQX4TH (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQXLTH (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQXLTH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRX1TH (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFRX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRX2TH (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFRX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRX4TH (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFRX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRXLTH (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFRXLTH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRHQX1TH (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFRHQX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRHQX2TH (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFRHQX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRHQX4TH (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFRHQX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRHQX8TH (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFRHQX8TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRQX1TH (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFRQX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRQX2TH (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFRQX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRQX4TH (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFRQX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRQXLTH (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN, tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN, tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFRQXLTH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSX1TH (Q, QN, D, SI, SE, CK, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

endspecify
endmodule // SDFFSX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSX2TH (Q, QN, D, SI, SE, CK, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

endspecify
endmodule // SDFFSX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSX4TH (Q, QN, D, SI, SE, CK, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

endspecify
endmodule // SDFFSX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSXLTH (Q, QN, D, SI, SE, CK, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

endspecify
endmodule // SDFFSXLTH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSHQX1TH (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSHQX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSHQX2TH (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSHQX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSHQX4TH (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSHQX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSHQX8TH (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSHQX8TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQX1TH (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSQX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQX2TH (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSQX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQX4TH (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSQX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQXLTH (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSQXLTH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRX1TH (Q, QN, D, SI, SE, CK, SN, RN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFSRX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRX2TH (Q, QN, D, SI, SE, CK, SN, RN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFSRX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRX4TH (Q, QN, D, SI, SE, CK, SN, RN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFSRX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRXLTH (Q, QN, D, SI, SE, CK, SN, RN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  not     N2 (QN, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN);

endspecify
endmodule // SDFFSRXLTH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX1TH (Q, D, SI, SE, CK, SN, RN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFSRHQX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX2TH (Q, D, SI, SE, CK, SN, RN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFSRHQX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX4TH (Q, D, SI, SE, CK, SN, RN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFSRHQX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX8TH (Q, D, SI, SE, CK, SN, RN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dSN;
wire dRN;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$RN$SN = 1.0,
      thold$SN$RN = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge RN &&& (SN == 1'b1), tsetup$RN$CK ,thold$RN$CK , NOTIFIER, , ,dCK,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER, , ,dCK,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(posedge RN, posedge SN, thold$SN$RN, NOTIFIER);    
    $hold(posedge SN, posedge RN, thold$RN$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q);

endspecify
endmodule // SDFFSRHQX8TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFTRX1TH (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);
   buf        I3 (scan, dSE);
   and        I4 (DandRN, dD, dRN);
   xor        I5 (flag, DandRN, dSI);
   not        I6 (notscan, dSE);
   and        I7 (checkD,dRN,notscan);
   and        I8 (scanD,dSI,dSE);
   and       I9 (DRN,dD,dRN);
   and        I10 (normD,DRN,notscan);
   or        I11 (Deff,scanD,normD);
   buf        I12 (checkRN,notscan);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
	(posedge CK *> (Q    +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
	(posedge CK *> (QN   -: Deff)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
     $setuphold(posedge CK &&& (checkD == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (checkD == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (checkRN == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (checkRN == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK, thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK, thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);

     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);


endspecify
endmodule // SDFFTRX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFTRX2TH (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);
   buf        I3 (scan, dSE);
   and        I4 (DandRN, dD, dRN);
   xor        I5 (flag, DandRN, dSI);
   not        I6 (notscan, dSE);
   and        I7 (checkD,dRN,notscan);
   and        I8 (scanD,dSI,dSE);
   and       I9 (DRN,dD,dRN);
   and        I10 (normD,DRN,notscan);
   or        I11 (Deff,scanD,normD);
   buf        I12 (checkRN,notscan);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
	(posedge CK *> (Q    +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
	(posedge CK *> (QN   -: Deff)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
     $setuphold(posedge CK &&& (checkD == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (checkD == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (checkRN == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (checkRN == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK, thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK, thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);

     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);


endspecify
endmodule // SDFFTRX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFTRX4TH (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);
   buf        I3 (scan, dSE);
   and        I4 (DandRN, dD, dRN);
   xor        I5 (flag, DandRN, dSI);
   not        I6 (notscan, dSE);
   and        I7 (checkD,dRN,notscan);
   and        I8 (scanD,dSI,dSE);
   and       I9 (DRN,dD,dRN);
   and        I10 (normD,DRN,notscan);
   or        I11 (Deff,scanD,normD);
   buf        I12 (checkRN,notscan);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
	(posedge CK *> (Q    +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
	(posedge CK *> (QN   -: Deff)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
     $setuphold(posedge CK &&& (checkD == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (checkD == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (checkRN == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (checkRN == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK, thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK, thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);

     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);


endspecify
endmodule // SDFFTRX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFTRXLTH (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
wire dRN;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);
   buf        I3 (scan, dSE);
   and        I4 (DandRN, dD, dRN);
   xor        I5 (flag, DandRN, dSI);
   not        I6 (notscan, dSE);
   and        I7 (checkD,dRN,notscan);
   and        I8 (scanD,dSI,dSE);
   and       I9 (DRN,dD,dRN);
   and        I10 (normD,DRN,notscan);
   or        I11 (Deff,scanD,normD);
   buf        I12 (checkRN,notscan);
  specify
    specparam 
      tplh$RN$Q = 1.0,
      tphl$RN$Q = 1.0,
      tplh$RN$QN = 1.0,
      tphl$RN$QN = 1.0,
      tminpwl$RN = 1.0,
      tminpwh$RN = 1.0,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
	(posedge CK *> (Q    +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
	(posedge CK *> (QN   -: Deff)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
     $setuphold(posedge CK &&& (checkD == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (checkD == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (checkRN == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (checkRN == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK, thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK, thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);

     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);


endspecify
endmodule // SDFFTRXLTH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFYQX2TH (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
wire dD;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_dff I0 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I1 (n1, dD, dSI, dSE);
  buf     I2 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, dD, dSI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFYQX2TH
`endcelldefine
	

//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFX1TH (Q, QN, D, CK, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);
  and     I3 (SandR, dSN, dRN);
  and     I4 (SandRandSE, SandR, dSE);
  not     I5 (SEb, dSE);
  and     I6 (SandRandSEbandE, SandR, SEb, dE);
  xor     I7 (DxorSI, dD, dSI);
  and     I8 (flag, DxorSI, SandR);
  and     I9 (SandRandSEb, SandR, SEb);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
    if (SandRandSEbandE == 1)
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (SandRandSE == 1)
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if (SandRandSEbandE == 1)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if (SandRandSE == 1)
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (SandRandSEbandE == 1), posedge D  , tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEbandE == 1), negedge D  , tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI ,  tsetup$SI$CK ,thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI ,  tsetup$SI$CK ,thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (flag == 1), posedge SE , tsetup$SE$CK , thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag == 1), negedge SE , tsetup$SE$CK , thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge E , tsetup$E$CK , thold$E$CK , NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge E ,  tsetup$E$CK ,thold$E$CK , NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFX1TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFX2TH (Q, QN, D, CK, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);
  and     I3 (SandR, dSN, dRN);
  and     I4 (SandRandSE, SandR, dSE);
  not     I5 (SEb, dSE);
  and     I6 (SandRandSEbandE, SandR, SEb, dE);
  xor     I7 (DxorSI, dD, dSI);
  and     I8 (flag, DxorSI, SandR);
  and     I9 (SandRandSEb, SandR, SEb);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
    if (SandRandSEbandE == 1)
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (SandRandSE == 1)
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if (SandRandSEbandE == 1)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if (SandRandSE == 1)
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (SandRandSEbandE == 1), posedge D  , tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEbandE == 1), negedge D  , tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI ,  tsetup$SI$CK ,thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI ,  tsetup$SI$CK ,thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (flag == 1), posedge SE , tsetup$SE$CK , thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag == 1), negedge SE , tsetup$SE$CK , thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge E , tsetup$E$CK , thold$E$CK , NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge E ,  tsetup$E$CK ,thold$E$CK , NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFX2TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFX4TH (Q, QN, D, CK, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);
  and     I3 (SandR, dSN, dRN);
  and     I4 (SandRandSE, SandR, dSE);
  not     I5 (SEb, dSE);
  and     I6 (SandRandSEbandE, SandR, SEb, dE);
  xor     I7 (DxorSI, dD, dSI);
  and     I8 (flag, DxorSI, SandR);
  and     I9 (SandRandSEb, SandR, SEb);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
    if (SandRandSEbandE == 1)
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (SandRandSE == 1)
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if (SandRandSEbandE == 1)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if (SandRandSE == 1)
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (SandRandSEbandE == 1), posedge D  , tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEbandE == 1), negedge D  , tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI ,  tsetup$SI$CK ,thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI ,  tsetup$SI$CK ,thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (flag == 1), posedge SE , tsetup$SE$CK , thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag == 1), negedge SE , tsetup$SE$CK , thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge E , tsetup$E$CK , thold$E$CK , NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge E ,  tsetup$E$CK ,thold$E$CK , NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFX4TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFXLTH (Q, QN, D, CK, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);
  and     I3 (SandR, dSN, dRN);
  and     I4 (SandRandSE, SandR, dSE);
  not     I5 (SEb, dSE);
  and     I6 (SandRandSEbandE, SandR, SEb, dE);
  xor     I7 (DxorSI, dD, dSI);
  and     I8 (flag, DxorSI, SandR);
  and     I9 (SandRandSEb, SandR, SEb);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
    if (SandRandSEbandE == 1)
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if (SandRandSE == 1)
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
    if (SandRandSEbandE == 1)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if (SandRandSE == 1)
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (SandRandSEbandE == 1), posedge D  , tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSEbandE == 1), negedge D  , tsetup$D$CK  ,thold$D$CK  , NOTIFIER, , ,dCK,dD);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI ,  tsetup$SI$CK ,thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI ,  tsetup$SI$CK ,thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (flag == 1), posedge SE , tsetup$SE$CK , thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag == 1), negedge SE , tsetup$SE$CK , thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge E , tsetup$E$CK , thold$E$CK , NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge E ,  tsetup$E$CK ,thold$E$CK , NOTIFIER, , ,dCK,dE);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFXLTH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFHQX1TH (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf       I1 (Q, n0);
   and       I3 (SandR, dSN, dRN);
   buf       I4 (scan, dSE);
   not       I5 (notscan, dSE);
   and       I6 (Dcheck, notscan, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
     if (notscan)
	(posedge CK *> (Q    +: E)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
	(posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     (posedge CK *> (Q    +: SE)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFHQX1TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFHQX2TH (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf       I1 (Q, n0);
   and       I3 (SandR, dSN, dRN);
   buf       I4 (scan, dSE);
   not       I5 (notscan, dSE);
   and       I6 (Dcheck, notscan, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
     if (notscan)
	(posedge CK *> (Q    +: E)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
	(posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     (posedge CK *> (Q    +: SE)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFHQX2TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFHQX4TH (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf       I1 (Q, n0);
   and       I3 (SandR, dSN, dRN);
   buf       I4 (scan, dSE);
   not       I5 (notscan, dSE);
   and       I6 (Dcheck, notscan, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
     if (notscan)
	(posedge CK *> (Q    +: E)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
	(posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     (posedge CK *> (Q    +: SE)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFHQX4TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFHQX8TH (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf       I1 (Q, n0);
   and       I3 (SandR, dSN, dRN);
   buf       I4 (scan, dSE);
   not       I5 (notscan, dSE);
   and       I6 (Dcheck, notscan, dE);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
     if (notscan)
	(posedge CK *> (Q    +: E)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
	(posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     (posedge CK *> (Q    +: SE)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFHQX8TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFTRX1TH (Q, QN, D, CK, E, SE, SI, RN);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);
   buf        I3 (scan, dSE);
   and        I4 (DandRN, dD, dRN);
   xor        I5 (flag, DandRN, dSI);
   not        I6 (notscan, dSE);
   and        I7 (Dcheck,dE,dRN,notscan);
   and        I8 (scanD,dSI,dSE);
   nand       I9 (DRN,dD,dRN);
   and        I10 (normD,DRN,notscan);
   nor        I11 (Deff,scanD,normD);
   buf        I15 (RNcheck, notscan);
   and        I14 (Echeck,dRN,notscan);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     (posedge CK *> (Q    +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
     (posedge CK *> (QN   -: Deff)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (Echeck == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (Echeck == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (RNcheck == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (RNcheck == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFTRX1TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFTRX2TH (Q, QN, D, CK, E, SE, SI, RN);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);
   buf        I3 (scan, dSE);
   and        I4 (DandRN, dD, dRN);
   xor        I5 (flag, DandRN, dSI);
   not        I6 (notscan, dSE);
   and        I7 (Dcheck,dE,dRN,notscan);
   and        I8 (scanD,dSI,dSE);
   nand       I9 (DRN,dD,dRN);
   and        I10 (normD,DRN,notscan);
   nor        I11 (Deff,scanD,normD);
   buf        I15 (RNcheck, notscan);
   and        I14 (Echeck,dRN,notscan);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     (posedge CK *> (Q    +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
     (posedge CK *> (QN   -: Deff)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (Echeck == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (Echeck == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (RNcheck == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (RNcheck == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFTRX2TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFTRX4TH (Q, QN, D, CK, E, SE, SI, RN);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);
   buf        I3 (scan, dSE);
   and        I4 (DandRN, dD, dRN);
   xor        I5 (flag, DandRN, dSI);
   not        I6 (notscan, dSE);
   and        I7 (Dcheck,dE,dRN,notscan);
   and        I8 (scanD,dSI,dSE);
   nand       I9 (DRN,dD,dRN);
   and        I10 (normD,DRN,notscan);
   nor        I11 (Deff,scanD,normD);
   buf        I15 (RNcheck, notscan);
   and        I14 (Echeck,dRN,notscan);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     (posedge CK *> (Q    +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
     (posedge CK *> (QN   -: Deff)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (Echeck == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (Echeck == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (RNcheck == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (RNcheck == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFTRX4TH
`endcelldefine


//$Id: edff.genpp,v 1.10 2006/03/27 16:02:32 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SEDFFTRXLTH (Q, QN, D, CK, E, SE, SI, RN);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
wire dD;
wire dCK;
wire dE;
wire dSE;
wire dSI;
wire dRN;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, dD, dCK, dRN, dSI, dSE, dE, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);
   buf        I3 (scan, dSE);
   and        I4 (DandRN, dD, dRN);
   xor        I5 (flag, DandRN, dSI);
   not        I6 (notscan, dSE);
   and        I7 (Dcheck,dE,dRN,notscan);
   and        I8 (scanD,dSI,dSE);
   nand       I9 (DRN,dD,dRN);
   and        I10 (normD,DRN,notscan);
   nor        I11 (Deff,scanD,normD);
   buf        I15 (RNcheck, notscan);
   and        I14 (Echeck,dRN,notscan);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      tsetup$RN$CK = 1.0,
      thold$RN$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     (posedge CK *> (Q    +: Deff)) = (tplh$CK$Q,  tphl$CK$Q);
     (posedge CK *> (QN   -: Deff)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER, , ,dCK,dD);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER, , ,dCK,dSI);
     $setuphold(posedge CK &&& (Echeck == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (Echeck == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
     $setuphold(posedge CK &&& (RNcheck == 1), posedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK &&& (RNcheck == 1), negedge RN, tsetup$RN$CK, thold$RN$CK, NOTIFIER, , ,dCK,dRN);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER, , ,dCK,dSE);
     $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK, tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK, tperiod$CK, NOTIFIER);
  endspecify
endmodule // SEDFFTRXLTH
`endcelldefine


//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SMDFFHQX1TH (Q, D0, D1, S0, SI, SE, CK);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff I1 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, dSI);
  xor     I12 (D0xorD1, dD0, dD1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (Q    +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb1 )
      (posedge CK *> (Q    +: D1)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER, , ,dCK,dS0);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER, , ,dCK,dS0);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SMDFFHQX1TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SMDFFHQX2TH (Q, D0, D1, S0, SI, SE, CK);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff I1 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, dSI);
  xor     I12 (D0xorD1, dD0, dD1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (Q    +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb1 )
      (posedge CK *> (Q    +: D1)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER, , ,dCK,dS0);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER, , ,dCK,dS0);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SMDFFHQX2TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SMDFFHQX4TH (Q, D0, D1, S0, SI, SE, CK);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff I1 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, dSI);
  xor     I12 (D0xorD1, dD0, dD1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (Q    +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb1 )
      (posedge CK *> (Q    +: D1)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER, , ,dCK,dS0);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER, , ,dCK,dS0);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SMDFFHQX4TH
`endcelldefine
	

//$Id: sdff.genpp,v 1.13 2006/03/27 16:02:02 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SMDFFHQX8TH (Q, D0, D1, S0, SI, SE, CK);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
wire dD0;
wire dD1;
wire dS0;
wire dSI;
wire dSE;
wire dCK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, dCK);
  udp_mux I0 (nm, dD0, dD1, dS0);
  udp_dff I1 (n0, n1, clk, dRN, dSN, NOTIFIER);
  udp_mux I2 (n1, nm, dSI, dSE);
  buf     I3 (Q, n0);
  and     I4 (SandR, dSN, dRN);
  and     I5 (SandRandSE, SandR, dSE);
  not     I6 (SEb, dSE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, dSI);
  xor     I12 (D0xorD1, dD0, dD1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (Q    +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb1 )
      (posedge CK *> (Q    +: D1)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER, , ,dCK,dD0);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER, , ,dCK,dD1);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER, , ,dCK,dSI);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER, , ,dCK,dS0);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER, , ,dCK,dS0);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SMDFFHQX8TH
`endcelldefine
	

//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TBUFX12TH (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // TBUFX12TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TBUFX16TH (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // TBUFX16TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TBUFX1TH (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // TBUFX1TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TBUFX20TH (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // TBUFX20TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TBUFX2TH (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // TBUFX2TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TBUFX3TH (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // TBUFX3TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TBUFX4TH (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // TBUFX4TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TBUFX6TH (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // TBUFX6TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TBUFX8TH (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // TBUFX8TH
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TBUFXLTH (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // TBUFXLTH
`endcelldefine
//$Id: tie.genpp,v 1.1.1.1 2002/12/05 17:56:00 ron Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TIEHITH (Y);
output Y;

  buf I0(Y, 1'b1);

endmodule //TIEHITH 
`endcelldefine
//$Id: tie.genpp,v 1.1.1.1 2002/12/05 17:56:00 ron Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TIELOTH (Y);
output Y;

  buf I0(Y, 1'b0);

endmodule //TIELOTH 
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATX1TH (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
wire dD;
wire dG;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not I3(clk,dG);
buf I4(flgclk,dG);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandR)
      (posedge G *> (QN -: D)) = (tplh$G$QN, tphl$G$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );

    // timing checks 5
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);


   endspecify
endmodule //TLATX1TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATX2TH (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
wire dD;
wire dG;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not I3(clk,dG);
buf I4(flgclk,dG);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandR)
      (posedge G *> (QN -: D)) = (tplh$G$QN, tphl$G$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );

    // timing checks 5
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);


   endspecify
endmodule //TLATX2TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATX4TH (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
wire dD;
wire dG;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not I3(clk,dG);
buf I4(flgclk,dG);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandR)
      (posedge G *> (QN -: D)) = (tplh$G$QN, tphl$G$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );

    // timing checks 5
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);


   endspecify
endmodule //TLATX4TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATXLTH (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
wire dD;
wire dG;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not I3(clk,dG);
buf I4(flgclk,dG);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandR)
      (posedge G *> (QN -: D)) = (tplh$G$QN, tphl$G$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );

    // timing checks 5
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);


   endspecify
endmodule //TLATXLTH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNX1TH (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
wire dD;
wire dGN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandR)
      (negedge GN *> (QN -: D)) = (tplh$GN$QN, tphl$GN$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );

    // timing checks 3
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);


   endspecify
endmodule //TLATNX1TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNX2TH (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
wire dD;
wire dGN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandR)
      (negedge GN *> (QN -: D)) = (tplh$GN$QN, tphl$GN$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );

    // timing checks 3
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);


   endspecify
endmodule //TLATNX2TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNX4TH (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
wire dD;
wire dGN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandR)
      (negedge GN *> (QN -: D)) = (tplh$GN$QN, tphl$GN$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );

    // timing checks 3
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);


   endspecify
endmodule //TLATNX4TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNXLTH (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
wire dD;
wire dGN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandR)
      (negedge GN *> (QN -: D)) = (tplh$GN$QN, tphl$GN$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );

    // timing checks 3
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);


   endspecify
endmodule //TLATNXLTH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNCAX12TH (ECK, E, CK);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK, posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //TLATNCAX12TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNCAX16TH (ECK, E, CK);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK, posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //TLATNCAX16TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNCAX20TH (ECK, E, CK);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK, posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //TLATNCAX20TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNCAX2TH (ECK, E, CK);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK, posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //TLATNCAX2TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNCAX3TH (ECK, E, CK);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK, posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //TLATNCAX3TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNCAX4TH (ECK, E, CK);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK, posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //TLATNCAX4TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNCAX6TH (ECK, E, CK);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK, posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //TLATNCAX6TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNCAX8TH (ECK, E, CK);
output ECK;
input  E, CK;
reg NOTIFIER;
wire dE;
wire dCK;

supply1 R, S;

  udp_tlat I0 (n0, dE, dCK, R, S, NOTIFIER);
  and      I1 (ECK, n0, CK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK, posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK, negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //TLATNCAX8TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNSRX1TH (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;
wire dD;
wire dGN;
wire dRN;
wire dSN;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tplh$RN$QN   = 1.0,
      tphl$RN$QN   = 1.0,
      tplh$SN$Q   = 1.0,
      tphl$SN$Q   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$GN$RN = 1.0,
      thold$GN$RN  = 0.5,
      tsetup$GN$SN = 1.0,
      thold$GN$SN  = 0.5,
      tsetup$RN$GN = 1.0,
      thold$RN$GN  = 0.5,
      tsetup$RN$SN = 1.0,
      thold$RN$SN  = 0.5,
      tsetup$SN$GN = 1.0,
      thold$SN$GN  = 0.5,
      tsetup$SN$RN = 1.0,
      thold$SN$RN  = 0.5,
      tminpwl$SN    = 1.0,
      tminpwl$RN    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandR)
      (negedge GN *> (QN -: D)) = (tplh$GN$QN, tphl$GN$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, posedge SN, tsetup$SN$GN,thold$SN$GN, NOTIFIER, , ,dGN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge GN, posedge RN &&& (SN == 1'b1), tsetup$RN$GN,thold$RN$GN, NOTIFIER, , ,dGN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 3
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    $hold(posedge RN, posedge SN, thold$SN$RN,NOTIFIER);
    $hold(posedge SN, posedge RN, thold$RN$SN,NOTIFIER);
    if (D == 1'b0 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && GN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && GN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && GN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && GN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule //TLATNSRX1TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNSRX2TH (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;
wire dD;
wire dGN;
wire dRN;
wire dSN;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tplh$RN$QN   = 1.0,
      tphl$RN$QN   = 1.0,
      tplh$SN$Q   = 1.0,
      tphl$SN$Q   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$GN$RN = 1.0,
      thold$GN$RN  = 0.5,
      tsetup$GN$SN = 1.0,
      thold$GN$SN  = 0.5,
      tsetup$RN$GN = 1.0,
      thold$RN$GN  = 0.5,
      tsetup$RN$SN = 1.0,
      thold$RN$SN  = 0.5,
      tsetup$SN$GN = 1.0,
      thold$SN$GN  = 0.5,
      tsetup$SN$RN = 1.0,
      thold$SN$RN  = 0.5,
      tminpwl$SN    = 1.0,
      tminpwl$RN    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandR)
      (negedge GN *> (QN -: D)) = (tplh$GN$QN, tphl$GN$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, posedge SN, tsetup$SN$GN,thold$SN$GN, NOTIFIER, , ,dGN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge GN, posedge RN &&& (SN == 1'b1), tsetup$RN$GN,thold$RN$GN, NOTIFIER, , ,dGN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 3
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    $hold(posedge RN, posedge SN, thold$SN$RN,NOTIFIER);
    $hold(posedge SN, posedge RN, thold$RN$SN,NOTIFIER);
    if (D == 1'b0 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && GN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && GN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && GN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && GN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule //TLATNSRX2TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNSRX4TH (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;
wire dD;
wire dGN;
wire dRN;
wire dSN;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tplh$RN$QN   = 1.0,
      tphl$RN$QN   = 1.0,
      tplh$SN$Q   = 1.0,
      tphl$SN$Q   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$GN$RN = 1.0,
      thold$GN$RN  = 0.5,
      tsetup$GN$SN = 1.0,
      thold$GN$SN  = 0.5,
      tsetup$RN$GN = 1.0,
      thold$RN$GN  = 0.5,
      tsetup$RN$SN = 1.0,
      thold$RN$SN  = 0.5,
      tsetup$SN$GN = 1.0,
      thold$SN$GN  = 0.5,
      tsetup$SN$RN = 1.0,
      thold$SN$RN  = 0.5,
      tminpwl$SN    = 1.0,
      tminpwl$RN    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandR)
      (negedge GN *> (QN -: D)) = (tplh$GN$QN, tphl$GN$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, posedge SN, tsetup$SN$GN,thold$SN$GN, NOTIFIER, , ,dGN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge GN, posedge RN &&& (SN == 1'b1), tsetup$RN$GN,thold$RN$GN, NOTIFIER, , ,dGN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 3
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    $hold(posedge RN, posedge SN, thold$SN$RN,NOTIFIER);
    $hold(posedge SN, posedge RN, thold$RN$SN,NOTIFIER);
    if (D == 1'b0 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && GN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && GN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && GN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && GN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule //TLATNSRX4TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNSRXLTH (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;
wire dD;
wire dGN;
wire dRN;
wire dSN;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, dGN);
not      I4 (flgclk, dGN);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tplh$RN$QN   = 1.0,
      tphl$RN$QN   = 1.0,
      tplh$SN$Q   = 1.0,
      tphl$SN$Q   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$GN$RN = 1.0,
      thold$GN$RN  = 0.5,
      tsetup$GN$SN = 1.0,
      thold$GN$SN  = 0.5,
      tsetup$RN$GN = 1.0,
      thold$RN$GN  = 0.5,
      tsetup$RN$SN = 1.0,
      thold$RN$SN  = 0.5,
      tsetup$SN$GN = 1.0,
      thold$SN$GN  = 0.5,
      tsetup$SN$RN = 1.0,
      thold$SN$RN  = 0.5,
      tminpwl$SN    = 1.0,
      tminpwl$RN    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandR)
      (negedge GN *> (QN -: D)) = (tplh$GN$QN, tphl$GN$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, posedge SN, tsetup$SN$GN,thold$SN$GN, NOTIFIER, , ,dGN,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge GN, posedge RN &&& (SN == 1'b1), tsetup$RN$GN,thold$RN$GN, NOTIFIER, , ,dGN,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 3
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER, , ,dGN,dD);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    $hold(posedge RN, posedge SN, thold$SN$RN,NOTIFIER);
    $hold(posedge SN, posedge RN, thold$RN$SN,NOTIFIER);
    if (D == 1'b0 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && GN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && GN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && GN == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && GN == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && GN == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && GN == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule //TLATNSRXLTH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNTSCAX12TH (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
  endspecify

endmodule //TLATNTSCAX12TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNTSCAX16TH (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
  endspecify

endmodule //TLATNTSCAX16TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNTSCAX20TH (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
  endspecify

endmodule //TLATNTSCAX20TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNTSCAX2TH (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
  endspecify

endmodule //TLATNTSCAX2TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNTSCAX3TH (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
  endspecify

endmodule //TLATNTSCAX3TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNTSCAX4TH (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
  endspecify

endmodule //TLATNTSCAX4TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNTSCAX6TH (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
  endspecify

endmodule //TLATNTSCAX6TH
`endcelldefine
//$Id: ckgate.genpp,v 1.9 2006/03/24 11:24:11 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATNTSCAX8TH (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;
wire dE;
wire dSE;
wire dCK;

supply1 R, S;

  or       I0 (n1, dSE, dE);
  udp_tlat I1 (n0, n1, dCK, R, S, NOTIFIER);
  and      I2 (ECK, n0, dCK);

  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      (posedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);
      (negedge CK *> (ECK  +: E)) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER, , ,dCK,dE);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER, , ,dCK,dSE);
  endspecify

endmodule //TLATNTSCAX8TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATSRX1TH (Q, QN, D, G, SN, RN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;
wire dD;
wire dG;
wire dSN;
wire dRN;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not I3(clk,dG);
buf I4(flgclk,dG);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$SN$Q   = 1.0,
      tphl$SN$Q   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tplh$RN$QN   = 1.0,
      tphl$RN$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$G$SN = 1.0,
      thold$G$SN  = 0.5,
      tsetup$G$RN = 1.0,
      thold$G$RN  = 0.5,
      tsetup$SN$G = 1.0,
      thold$SN$G  = 0.5,
      tsetup$SN$RN = 1.0,
      thold$SN$RN  = 0.5,
      tsetup$RN$G = 1.0,
      thold$RN$G  = 0.5,
      tsetup$RN$SN = 1.0,
      thold$RN$SN  = 0.5,
      tminpwl$SN    = 1.0,
      tminpwl$RN    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandR)
      (posedge G *> (QN -: D)) = (tplh$G$QN, tphl$G$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, posedge SN, tsetup$SN$G,thold$SN$G, NOTIFIER, , ,dG,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge G, posedge RN &&& (SN == 1'b1), tsetup$RN$G,thold$RN$G, NOTIFIER, , ,dG,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 5
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

    $hold(posedge RN, posedge SN, thold$SN$RN,NOTIFIER);
    $hold(posedge SN, posedge RN, thold$RN$SN,NOTIFIER);
    if (D == 1'b0 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && G == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && G == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && G == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && G == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule //TLATSRX1TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATSRX2TH (Q, QN, D, G, SN, RN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;
wire dD;
wire dG;
wire dSN;
wire dRN;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not I3(clk,dG);
buf I4(flgclk,dG);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$SN$Q   = 1.0,
      tphl$SN$Q   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tplh$RN$QN   = 1.0,
      tphl$RN$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$G$SN = 1.0,
      thold$G$SN  = 0.5,
      tsetup$G$RN = 1.0,
      thold$G$RN  = 0.5,
      tsetup$SN$G = 1.0,
      thold$SN$G  = 0.5,
      tsetup$SN$RN = 1.0,
      thold$SN$RN  = 0.5,
      tsetup$RN$G = 1.0,
      thold$RN$G  = 0.5,
      tsetup$RN$SN = 1.0,
      thold$RN$SN  = 0.5,
      tminpwl$SN    = 1.0,
      tminpwl$RN    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandR)
      (posedge G *> (QN -: D)) = (tplh$G$QN, tphl$G$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, posedge SN, tsetup$SN$G,thold$SN$G, NOTIFIER, , ,dG,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge G, posedge RN &&& (SN == 1'b1), tsetup$RN$G,thold$RN$G, NOTIFIER, , ,dG,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 5
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

    $hold(posedge RN, posedge SN, thold$SN$RN,NOTIFIER);
    $hold(posedge SN, posedge RN, thold$RN$SN,NOTIFIER);
    if (D == 1'b0 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && G == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && G == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && G == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && G == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule //TLATSRX2TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATSRX4TH (Q, QN, D, G, SN, RN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;
wire dD;
wire dG;
wire dSN;
wire dRN;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not I3(clk,dG);
buf I4(flgclk,dG);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$SN$Q   = 1.0,
      tphl$SN$Q   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tplh$RN$QN   = 1.0,
      tphl$RN$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$G$SN = 1.0,
      thold$G$SN  = 0.5,
      tsetup$G$RN = 1.0,
      thold$G$RN  = 0.5,
      tsetup$SN$G = 1.0,
      thold$SN$G  = 0.5,
      tsetup$SN$RN = 1.0,
      thold$SN$RN  = 0.5,
      tsetup$RN$G = 1.0,
      thold$RN$G  = 0.5,
      tsetup$RN$SN = 1.0,
      thold$RN$SN  = 0.5,
      tminpwl$SN    = 1.0,
      tminpwl$RN    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandR)
      (posedge G *> (QN -: D)) = (tplh$G$QN, tphl$G$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, posedge SN, tsetup$SN$G,thold$SN$G, NOTIFIER, , ,dG,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge G, posedge RN &&& (SN == 1'b1), tsetup$RN$G,thold$RN$G, NOTIFIER, , ,dG,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 5
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

    $hold(posedge RN, posedge SN, thold$SN$RN,NOTIFIER);
    $hold(posedge SN, posedge RN, thold$RN$SN,NOTIFIER);
    if (D == 1'b0 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && G == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && G == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && G == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && G == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule //TLATSRX4TH
`endcelldefine
//$Id: tlat.genpp,v 1.8 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TLATSRXLTH (Q, QN, D, G, SN, RN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;
wire dD;
wire dG;
wire dSN;
wire dRN;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, dD, clk, dRN, dSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not I3(clk,dG);
buf I4(flgclk,dG);
and      I5 (SandR, dSN, dRN);
and      I6 (SandRandCLK, dSN,dRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$SN$Q   = 1.0,
      tphl$SN$Q   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tplh$RN$QN   = 1.0,
      tphl$RN$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$G$SN = 1.0,
      thold$G$SN  = 0.5,
      tsetup$G$RN = 1.0,
      thold$G$RN  = 0.5,
      tsetup$SN$G = 1.0,
      thold$SN$G  = 0.5,
      tsetup$SN$RN = 1.0,
      thold$SN$RN  = 0.5,
      tsetup$RN$G = 1.0,
      thold$RN$G  = 0.5,
      tsetup$RN$SN = 1.0,
      thold$RN$SN  = 0.5,
      tminpwl$SN    = 1.0,
      tminpwl$RN    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandR)
      (posedge G *> (QN -: D)) = (tplh$G$QN, tphl$G$QN);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, posedge SN, tsetup$SN$G,thold$SN$G, NOTIFIER, , ,dG,dSN);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge G, posedge RN &&& (SN == 1'b1), tsetup$RN$G,thold$RN$G, NOTIFIER, , ,dG,dRN);
    $width(negedge RN &&& (SN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 5
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER, , ,dG,dD);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

    $hold(posedge RN, posedge SN, thold$SN$RN,NOTIFIER);
    $hold(posedge SN, posedge RN, thold$RN$SN,NOTIFIER);
    if (D == 1'b0 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b1 && G == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (Q +: 1'b0)) = (tplh$RN$Q, tphl$RN$Q); 
    if (D == 1'b0 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && G == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && G == 1'b0 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b1 && G == 1'b1 && SN == 1'b1 )
       (negedge  RN *> (QN -: 1'b0)) = (tplh$RN$QN, tphl$RN$QN); 
    if (D == 1'b0 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b1 && G == 1'b0 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN); 
    if (D == 1'b0 && G == 1'b1 && RN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);

   endspecify
endmodule //TLATSRXLTH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2X1TH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2X1TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2X2TH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2X2TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2X4TH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2X4TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2XLTH (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2XLTH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3X1TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3X1TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3X2TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3X2TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3X4TH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3X4TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3XLTH (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3XLTH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X1TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X1TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X2TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X2TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X3TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X3TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X4TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X4TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X8TH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X8TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2XLTH (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2XLTH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3X1TH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3X1TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3X2TH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3X2TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3X4TH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3X4TH
`endcelldefine
//$Id: xor.genpp,v 1.4 2006/01/09 06:34:38 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3XLTH (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3XLTH
`endcelldefine


primitive udp_sedff (out, in, clk, clr_, si, se, en, NOTIFIER);
   output out;  
   input  in, clk, clr_, si, se,  en, NOTIFIER;
   reg    out;

   table
   // in  clk  clr_  si  se  en  NOT : Qt : Qt+1
      ?    ?    ?     ?   ?   ?   *  : ?  :  x; // any notifier changed
      ?    ?    0     ?   ?   ?   ?  : ?  :  0;     
      ?    r    ?     0   1   ?   ?  : ?  :  0;     
      ?    r    1     1   1   ?   ?  : ?  :  1;
      ?    b    1     ?   *   ?   ?  : ?  :  -; // no changes when se switches
      ?    b    1     *   ?   ?   ?  : ?  :  -; // no changes when si switches
      *    b    1     ?   ?   ?   ?  : ?  :  -; // no changes when in switches
      *    ?    ?     ?   0   0   ?  : 0  :  0; // no changes when in switches
      ?    ?    ?     *   0   0   ?  : 0  :  0; // no changes when in switches
      ?    b    1     ?   ?   *   ?  : ?  :  -; // no changes when en switches
      ?    b    *     ?   ?   ?   ?  : 0  :  0; // no changes when en switches
      ?    ?    *     ?   0   0   ?  : 0  :  0; // no changes when en switches
      ?    b    ?     ?   ?   *   ?  : 0  :  0; // no changes when en switches
      ?    b    ?     ?   *   ?   ?  : 0  :  0; // no changes when en switches
      ?    b    ?     *   ?   ?   ?  : 0  :  0; // no changes when en switches
      *    b    ?     ?   ?   ?   ?  : 0  :  0; // no changes when en switches
      ?  (10)   ?     ?   ?   ?   ?  : ?  :  -;  // no changes on falling clk edge
      ?    *    1     1   1   ?   ?  : 1  :  1;
      ?    x    1     1   1   ?   ?  : 1  :  1;
      ?    *    1     1   ?   0   ?  : 1  :  1;
      ?    x    1     1   ?   0   ?  : 1  :  1;
      ?    *    ?     0   1   ?   ?  : 0  :  0;
      ?    x    ?     0   1   ?   ?  : 0  :  0;
      ?    *    ?     0   ?   0   ?  : 0  :  0;
      ?    x    ?     0   ?   0   ?  : 0  :  0;
      0    r    ?     0   ?   1   ?  : ?  :  0 ; 
      0    *    ?     0   ?   ?   ?  : 0  :  0 ; 
      0    x    ?     0   ?   ?   ?  : 0  :  0 ; 
      1    r    1     1   ?   1   ?  : ?  :  1 ; 
      1    *    1     1   ?   ?   ?  : 1  :  1 ; 
      1    x    1     1   ?   ?   ?  : 1  :  1 ; 
      ?  (x0)   ?     ?   ?   ?   ?  : ?  :  -;  // no changes on falling clk edge
      1    r    1     ?   0   1   ?  : ?  :  1;
      0    r    ?     ?   0   1   ?  : ?  :  0;
      ?    *    ?     ?   0   0   ?  : ?  :  -;
      ?    x    1     ?   0   0   ?  : ?  :  -;
      1    x    1     ?   0   ?   ?  : 1  :  1; // no changes when in switches
      0    x    ?     ?   0   ?   ?  : 0  :  0; // no changes when in switches
      1    x    ?     ?   0   0   ?  : 0  :  0; // no changes when in switches
      1    *    1     ?   0   ?   ?  : 1  :  1; // reduce pessimism
      0    *    ?     ?   0   ?   ?  : 0  :  0; // reduce pessimism

   endtable
endprimitive  /* udp_sedff */
   


primitive udp_edfft (out, in, clk, clr_, set_, en, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, en, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  en  NOT  : Qt : Qt+1
//
   ?   r    0      1     ?   ?    : ?  :  0  ; // clock in 0
   0   r    ?      1     1   ?    : ?  :  0  ; // clock in 0
   ?   r    ?      0     ?   ?    : ?  :  1  ; // clock in 1
   1   r    1      ?     1   ?    : ?  :  1  ; // clock in 1
   ?   *    1      1     0   ?    : ?  :  -  ; // no changes, not enabled
   ?   *    ?      1     0   ?    : 0  :  0  ; // no changes, not enabled
   ?   *    1      ?     0   ?    : 1  :  1  ; // no changes, not enabled
   ?  (x0)  ?      ?     ?   ?    : ?  :  -  ; // no changes
   ?  (x1)  ?      0     ?   ?    : 1  :  1  ; // no changes
   1   *    1      ?     ?   ?    : 1  :  1  ; // reduce pessimism
   0   *    ?      1     ?   ?    : 0  :  0  ; // reduce pessimism
   ?   f    ?      ?     ?   ?    : ?  :  -  ; // no changes on negedge clk
   *   b    ?      ?     ?   ?    : ?  :  -  ; // no changes when in switches
   1   x    1      ?     ?   ?    : 1  :  1  ; // no changes when in switches
   ?   x    1      ?     0   ?    : 1  :  1  ; // no changes when in switches
   0   x    ?      1     ?   ?    : 0  :  0  ; // no changes when in switches
   ?   x    ?      1     0   ?    : 0  :  0  ; // no changes when in switches
   ?   b    ?      ?     *   ?    : ?  :  -  ; // no changes when en switches
   ?   b    *      ?     ?   ?    : ?  :  -  ; // no changes when clr_ switches
   ?   x    0      1     ?   ?    : 0  :  0  ; // no changes when clr_ switches
   ?   b    ?      *     ?   ?    : ?  :  -  ; // no changes when set_ switches
   ?   x    ?      0     ?   ?    : 1  :  1  ; // no changes when set_ switches
   ?   ?    ?      ?     ?   *    : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_edfft


primitive udp_mux (out, in, s_in, s_sel);
   output out;  
   input  in, s_in, s_sel;

   table

// in  s_in  s_sel :  out
//
   1  ?   0  :  1 ;
   0  ?   0  :  0 ;
   ?  1   1  :  1 ;
   ?  0   1  :  0 ;
   0  0   x  :  0 ;
   1  1   x  :  1 ;

   endtable
endprimitive // udp_mux


primitive udp_sedfft (out, in, clk, clr_, si, se, en, NOTIFIER);
   output out;  
   input  in, clk, clr_, si, se,  en, NOTIFIER;
   reg    out;

   table
   // in  clk  clr_  si  se  en  NOT : Qt : Qt+1
      ?    ?    ?     ?   ?   ?   *  : ?  :  x; // any notifier changed
      ?    r    ?     0   1   ?   ?  : ?  :  0;     
      ?    r    ?     1   1   ?   ?  : ?  :  1;
      ?    b    ?     ?   *   ?   ?  : ?  :  -; // no changes when se switches
      ?    b    ?     *   ?   ?   ?  : ?  :  -; // no changes when si switches
      *    b    ?     ?   ?   ?   ?  : ?  :  -; // no changes when in switches
      ?    b    ?     ?   ?   *   ?  : ?  :  -; // no changes when en switches
      ?    b    *     ?   ?   ?   ?  : ?  :  -; // no changes when clr switches
      0    r    ?     0   ?   1   ?  : ?  :  0 ; 
      1    r    1     1   ?   1   ?  : ?  :  1 ; 
      ?    r    ?     0   ?   0   ?  : 0  :  0;
      ?    x    ?     0   ?   0   ?  : 0  :  0;
      ?    r    1     1   ?   0   ?  : 1  :  1;
      ?    x    1     1   ?   0   ?  : 1  :  1;
      ?    *    1     ?   0   0   ?  : ?  :  -;
      ?    *    ?     1   1   ?   ?  : 1  :  1;
      1    *    1     1   ?   ?   ?  : 1  :  1;
      ?    *    ?     0   1   ?   ?  : 0  :  0;
      ?    *    0     0   ?   ?   ?  : 0  :  0;
      0    *    ?     0   ?   ?   ?  : 0  :  0;
      ?    x    1     ?   0   0   ?  : ?  :  -;
      ?    *    ?     ?   0   0   ?  : 0  :  0;
      ?    x    ?     ?   0   0   ?  : 0  :  0;
      ?    x    ?     1   1   ?   ?  : 1  :  1;
      1    x    1     1   ?   ?   ?  : 1  :  1;
      ?    x    ?     0   1   ?   ?  : 0  :  0;
      ?    x    0     0   ?   ?   ?  : 0  :  0;
      0    x    ?     0   ?   ?   ?  : 0  :  0;
      ?    r    0     0   ?   ?   ?  : ?  :  0 ; 
      ?   (?0)  ?     ?   ?   ?   ?  : ?  :  -;  // no changes on falling clk edge
      1    r    1     ?   0   1   ?  : ?  :  1;
      0    r    ?     ?   0   1   ?  : ?  :  0;
      ?    r    0     ?   0   ?   ?  : ?  :  0;
      ?    x    0     ?   0   ?   ?  : 0  :  0;
      1    x    1     ?   0   ?   ?  : 1  :  1; // no changes when in switches
      0    x    ?     ?   0   ?   ?  : 0  :  0; // no changes when in switches
      1    *    1     ?   0   ?   ?  : 1  :  1; // reduce pessimism
      0    *    ?     ?   0   ?   ?  : 0  :  0; // reduce pessimism

   endtable
endprimitive  /* udp_sedfft */
   


primitive udp_mux2 (out, in0, in1, sel);
   output out;  
   input  in0, in1, sel;

   table

// in0 in1  sel :  out
//
   1  ?   0  :  1 ;
   0  ?   0  :  0 ;
   ?  1   1  :  1 ;
   ?  0   1  :  0 ;
   0  0   x  :  0 ;
   1  1   x  :  1 ;

   endtable
endprimitive // udp_mux2


primitive udp_tlatrf (out, in, ww, wwn, NOTIFIER);
   output out;  
   input  in, ww, wwn, NOTIFIER;
   reg    out;

   table

// in  ww    wwn  NOT  : Qt : Qt+1
//	     
   1   ?     0    ?    : ?  :  1  ; // 
   1   1     ?    ?    : ?  :  1  ; // 
   0   ?     0    ?    : ?  :  0  ; // 
   0   1     ?    ?    : ?  :  0  ; // 
   1   *     ?    ?    : 1  :  1  ; // reduce pessimism
   1   ?     *    ?    : 1  :  1  ; // reduce pessimism
   0   *     ?    ?    : 0  :  0  ; // reduce pessimism
   0   ?     *    ?    : 0  :  0  ; // reduce pessimism
   *   0     1    ?    : ?  :  -  ; // no changes when in switches
   ?   ?     ?    *    : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_tlatrf



primitive udp_mux4 (out, in0, in1, in2, in3, sel_0, sel_1);
   output out;  
   input  in0, in1, in2, in3, sel_0, sel_1;

   table

// in0 in1 in2 in3 sel_0 sel_1 :  out
//
   0  ?  ?  ?  0  0  :  0;
   1  ?  ?  ?  0  0  :  1;
   ?  0  ?  ?  1  0  :  0;
   ?  1  ?  ?  1  0  :  1;
   ?  ?  0  ?  0  1  :  0;
   ?  ?  1  ?  0  1  :  1;
   ?  ?  ?  0  1  1  :  0;
   ?  ?  ?  1  1  1  :  1;
   0  0  ?  ?  x  0  :  0;
   1  1  ?  ?  x  0  :  1;
   ?  ?  0  0  x  1  :  0;
   ?  ?  1  1  x  1  :  1;
   0  ?  0  ?  0  x  :  0;
   1  ?  1  ?  0  x  :  1;
   ?  0  ?  0  1  x  :  0;
   ?  1  ?  1  1  x  :  1;
   1  1  1  1  x  x  :  1;
   0  0  0  0  x  x  :  0;

   endtable
endprimitive // udp_mux4


primitive udp_dff (out, in, clk, clr_, set_, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  NOT  : Qt : Qt+1
//
   0  r   ?   1   ?   : ?  :  0  ; // clock in 0
   1  r   1   ?   ?   : ?  :  1  ; // clock in 1
   1  *   1   ?   ?   : 1  :  1  ; // reduce pessimism
   0  *   ?   1   ?   : 0  :  0  ; // reduce pessimism
   ?  f   ?   ?   ?   : ?  :  -  ; // no changes on negedge clk
   *  b   ?   ?   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   ?   0   ?   : ?  :  1  ; // set output
   ?  b   1   *   ?   : 1  :  1  ; // cover all transistions on set_
   1  x   1   *   ?   : 1  :  1  ; // cover all transistions on set_
   ?  ?   0   1   ?   : ?  :  0  ; // reset output
   ?  b   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
   0  x   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_dff


primitive udp_outrf (out, in, rwn, rw);
   output out;  
   input  in, rwn, rw;

   table

// in  rwn   rw   : out;
//	     	  
   0   0     ?    : 1  ; // 
   1   ?     1    : 1  ; // 
   ?   1     0    : 0  ; // 
   1   ?     0    : 0  ; // 
   0   1     ?    : 0  ; // 

   endtable
endprimitive // udp_outrf



primitive udp_tlat (out, in, hold, clr_, set_, NOTIFIER);
   output out;  
   input  in, hold, clr_, set_, NOTIFIER;
   reg    out;

   table

// in  hold  clr_   set_  NOT  : Qt : Qt+1
//
   1  0   1   ?   ?   : ?  :  1  ; // 
   0  0   ?   1   ?   : ?  :  0  ; // 
   1  *   1   ?   ?   : 1  :  1  ; // reduce pessimism
   0  *   ?   1   ?   : 0  :  0  ; // reduce pessimism
   *  1   ?   ?   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   ?   0   ?   : ?  :  1  ; // set output
   ?  1   1   *   ?   : 1  :  1  ; // cover all transistions on set_
   1  ?   1   *   ?   : 1  :  1  ; // cover all transistions on set_
   ?  ?   0   1   ?   : ?  :  0  ; // reset output
   ?  1   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
   0  ?   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_tlat


primitive udp_edff (out, in, clk, clr_, set_, en, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, en, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  en  NOT  : Qt : Qt+1
//
   0   r    ?      1     1   ?    : ?  :  0  ; // clock in 0
   1   r    1      ?     1   ?    : ?  :  1  ; // clock in 1
   ?   *    ?      ?     0   ?    : ?  :  -  ; // no changes, not enabled
   *   ?    ?      ?     0   ?    : ?  :  -  ; // no changes, not enabled
   1   *    1      ?     ?   ?    : 1  :  1  ; // reduce pessimism
   0   *    ?      1     ?   ?    : 0  :  0  ; // reduce pessimism
   ?   f    ?      ?     ?   ?    : ?  :  -  ; // no changes on negedge clk
   *   b    ?      ?     ?   ?    : ?  :  -  ; // no changes when in switches
   1   x    1      ?     ?   ?    : 1  :  1  ; // no changes when in switches
   0   x    ?      1     ?   ?    : 0  :  0  ; // no changes when in switches
   ?   b    ?      ?     *   ?    : ?  :  -  ; // no changes when en switches
   ?   x    1      1     0   ?    : ?  :  -  ; // no changes when en is disabled
   ?   ?    ?      0     ?   ?    : ?  :  1  ; // set output
   ?   b    1      *     ?   ?    : 1  :  1  ; // cover all transistions on set_
   ?   ?    1      *     0   ?    : 1  :  1  ; // cover all transistions on set_
   ?   ?    0      1     ?   ?    : ?  :  0  ; // reset output
   ?   b    *      1     ?   ?    : 0  :  0  ; // cover all transistions on clr_
   ?   ?    *      1     0   ?    : 0  :  0  ; // cover all transistions on clr_
   ?   ?    ?      ?     ?   *    : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_edff


primitive udp_bmx (out, x2, a, s, m1, m0);
   output out;  
   input   x2, a, s, m1, m0;

   table

// x2 a  s m1 m0 :  out
//
   0  1  0  0  ? :  1;
   0  1  0  1  ? :  0;
   0  0  1  0  ? :  0;
   0  0  1  1  ? :  1;
   1  1  0  ?  0 :  1;
   1  1  0  ?  1 :  0;
   1  0  1  ?  0 :  0;
   1  0  1  ?  1 :  1;
   ?  0  0  ?  ? :  1;
   ?  1  1  ?  ? :  0;
   ?  ?  1  0  0 :  0;
   ?  0  ?  1  1 :  1;
   ?  ?  0  0  0 :  1;
   ?  1  ?  1  1 :  0;

   endtable
endprimitive // udp_bmx
